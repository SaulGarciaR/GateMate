//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (28 Feb 2023)
//  Compile Time: 2023-02-28 18:50:27
//  Program Run:  2023-08-04 13:33:24
//  Program Call: ../../bin/p_r/p_r -i net/aes256_uart_synth.v -o aes256_uart -ccf src/aes256_uart.ccf 
//  File Type:    Verilog

// Gatecount:   3696
module aes256_uart (clk , data_in , reset_n ,
       data_out , led 
       ) ;

input  clk;
input  data_in;
input  reset_n;

output data_out;
output [5:0]led;



wire [5:0]led;
wire clk;
wire data_in;
wire na1_1;
wire na2_1;
wire na3_2;
wire na4_1;
wire na5_2;
wire na6_1;
wire na7_2;
wire na8_1;
wire na9_2;
wire na10_1;
wire na11_2;
wire na12_1;
wire na13_1;
wire na14_1;
wire na15_2;
wire na16_2;
wire na17_1;
wire na18_1;
wire na19_1;
wire na20_1;
wire na21_2;
wire na22_2;
wire na23_1;
wire na24_2;
wire na25_1;
wire na26_2;
wire na27_1;
wire na28_1;
wire na30_1;
wire na31_1;
wire na32_2;
wire na33_1;
wire na34_1;
wire na36_1;
wire na37_1;
wire na38_1;
wire na39_1;
wire na40_1;
wire na42_1;
wire na43_1;
wire na44_2;
wire na45_1;
wire na46_1;
wire na48_1;
wire na49_1;
wire na50_1;
wire na51_1;
wire na52_1;
wire na54_1;
wire na55_1;
wire na56_2;
wire na57_2;
wire na58_1;
wire na59_1;
wire na61_1;
wire na62_1;
wire na63_2;
wire na64_1;
wire na65_1;
wire na67_1;
wire na68_1;
wire na69_1;
wire na70_1;
wire na71_1;
wire na73_2;
wire na74_1;
wire na75_1;
wire na76_1;
wire na77_1;
wire na79_2;
wire na80_1;
wire na81_1;
wire na82_1;
wire na83_1;
wire na85_1;
wire na86_1;
wire na87_1;
wire na88_1;
wire na89_1;
wire na91_1;
wire na92_1;
wire na93_1;
wire na94_1;
wire na95_1;
wire na97_1;
wire na98_1;
wire na99_1;
wire na100_1;
wire na101_1;
wire na103_1;
wire na105_1;
wire na106_1;
wire na107_1;
wire na109_1;
wire na110_1;
wire na111_2;
wire na112_1;
wire na113_1;
wire na115_2;
wire na116_1;
wire na117_1;
wire na118_1;
wire na119_1;
wire na121_2;
wire na122_1;
wire na123_1;
wire na124_1;
wire na125_1;
wire na127_1;
wire na128_1;
wire na129_1;
wire na130_1;
wire na131_1;
wire na133_1;
wire na134_1;
wire na135_1;
wire na136_1;
wire na137_1;
wire na139_1;
wire na140_1;
wire na141_1;
wire na142_1;
wire na143_1;
wire na145_2;
wire na146_1;
wire na147_1;
wire na148_1;
wire na149_1;
wire na151_2;
wire na152_1;
wire na153_1;
wire na154_1;
wire na155_1;
wire na157_1;
wire na158_1;
wire na159_2;
wire na160_1;
wire na161_1;
wire na163_1;
wire na165_1;
wire na166_1;
wire na167_1;
wire na169_1;
wire na170_1;
wire na171_1;
wire na172_1;
wire na173_1;
wire na175_1;
wire na176_1;
wire na177_1;
wire na178_1;
wire na179_1;
wire na181_1;
wire na182_1;
wire na183_1;
wire na184_1;
wire na185_1;
wire na187_1;
wire na188_1;
wire na189_2;
wire na190_1;
wire na191_1;
wire na193_2;
wire na194_1;
wire na195_1;
wire na196_1;
wire na197_1;
wire na199_1;
wire na200_1;
wire na201_2;
wire na202_1;
wire na203_1;
wire na205_1;
wire na206_1;
wire na207_1;
wire na208_1;
wire na209_1;
wire na211_1;
wire na212_1;
wire na213_1;
wire na214_1;
wire na215_2;
wire na216_2;
wire na217_1;
wire na218_1;
wire na219_1;
wire na220_2;
wire na221_2;
wire na222_2;
wire na223_1;
wire na224_1;
wire na225_1;
wire na226_1;
wire na227_1;
wire na228_2;
wire na229_1;
wire na230_2;
wire na231_2;
wire na232_1;
wire na234_1;
wire na236_1;
wire na237_1;
wire na238_1;
wire na239_1;
wire na240_2;
wire na241_1;
wire na242_2;
wire na243_1;
wire na244_1;
wire na245_1;
wire na246_1;
wire na247_2;
wire na248_1;
wire na249_1;
wire na250_1;
wire na251_1;
wire na252_1;
wire na253_2;
wire na254_1;
wire na255_2;
wire na256_1;
wire na258_1;
wire na259_1;
wire na260_1;
wire na261_1;
wire na262_2;
wire na263_1;
wire na264_1;
wire na266_1;
wire na267_1;
wire na268_1;
wire na269_1;
wire na270_1;
wire na272_1;
wire na273_1;
wire na274_2;
wire na275_1;
wire na276_1;
wire na278_1;
wire na279_1;
wire na280_1;
wire na281_1;
wire na283_1;
wire na284_1;
wire na285_1;
wire na286_1;
wire na287_1;
wire na288_1;
wire na290_1;
wire na292_1;
wire na293_1;
wire na294_1;
wire na295_2;
wire na296_1;
wire na297_2;
wire na298_1;
wire na300_1;
wire na301_1;
wire na302_1;
wire na303_2;
wire na305_1;
wire na307_1;
wire na308_1;
wire na309_1;
wire na310_1;
wire na311_1;
wire na312_1;
wire na313_2;
wire na314_1;
wire na315_1;
wire na316_1;
wire na317_1;
wire na319_1;
wire na320_1;
wire na322_1;
wire na323_2;
wire na324_1;
wire na327_1;
wire na328_1;
wire na332_1;
wire na334_1;
wire na335_1;
wire na336_1;
wire na339_1;
wire na343_1;
wire na344_1;
wire na345_1;
wire na348_1;
wire na352_1;
wire na353_1;
wire na354_1;
wire na355_1;
wire na357_1;
wire na358_1;
wire na360_1;
wire na363_1;
wire na366_1;
wire na370_1;
wire na371_1;
wire na372_1;
wire na373_1;
wire na375_1;
wire na376_1;
wire na378_1;
wire na381_1;
wire na382_1;
wire na384_1;
wire na385_1;
wire na386_2;
wire na387_1;
wire na390_1;
wire na391_1;
wire na393_1;
wire na394_1;
wire na398_1;
wire na399_1;
wire na401_1;
wire na402_1;
wire na403_1;
wire na404_1;
wire na407_1;
wire na408_1;
wire na410_1;
wire na411_1;
wire na413_1;
wire na416_1;
wire na417_1;
wire na420_1;
wire na421_1;
wire na422_1;
wire na425_1;
wire na426_1;
wire na428_1;
wire na429_1;
wire na431_1;
wire na434_1;
wire na435_1;
wire na437_1;
wire na438_1;
wire na442_1;
wire na443_1;
wire na446_1;
wire na447_1;
wire na448_1;
wire na451_1;
wire na452_1;
wire na454_1;
wire na455_1;
wire na456_1;
wire na457_1;
wire na460_1;
wire na463_1;
wire na467_1;
wire na468_1;
wire na469_1;
wire na470_1;
wire na473_1;
wire na474_1;
wire na477_1;
wire na480_1;
wire na484_1;
wire na485_1;
wire na486_1;
wire na487_1;
wire na491_1;
wire na493_1;
wire na494_1;
wire na495_1;
wire na496_1;
wire na498_1;
wire na499_1;
wire na501_1;
wire na504_1;
wire na508_1;
wire na509_1;
wire na510_1;
wire na513_1;
wire na516_1;
wire na520_1;
wire na521_1;
wire na522_1;
wire na523_1;
wire na525_1;
wire na526_1;
wire na527_1;
wire na528_1;
wire na531_2;
wire na532_1;
wire na533_1;
wire na534_2;
wire na535_2;
wire na536_2;
wire na537_1;
wire na538_1;
wire na539_2;
wire na540_1;
wire na541_1;
wire na542_1;
wire na543_2;
wire na544_1;
wire na545_1;
wire na546_1;
wire na547_1;
wire na548_1;
wire na549_1;
wire na550_1;
wire na551_1;
wire na552_1;
wire na553_1;
wire na554_1;
wire na555_1;
wire na556_1;
wire na557_1;
wire na558_1;
wire na559_1;
wire na560_1;
wire na561_1;
wire na562_1;
wire na563_1;
wire na564_1;
wire na565_1;
wire na566_1;
wire na567_1;
wire na568_1;
wire na569_1;
wire na570_1;
wire na571_1;
wire na572_1;
wire na573_1;
wire na574_1;
wire na575_1;
wire na576_1;
wire na577_1;
wire na578_1;
wire na579_1;
wire na580_1;
wire na581_1;
wire na582_1;
wire na583_1;
wire na584_1;
wire na585_1;
wire na586_1;
wire na587_1;
wire na588_1;
wire na589_1;
wire na590_1;
wire na591_1;
wire na592_1;
wire na593_1;
wire na594_1;
wire na595_1;
wire na596_1;
wire na597_1;
wire na598_1;
wire na599_1;
wire na600_1;
wire na601_1;
wire na602_1;
wire na603_1;
wire na604_1;
wire na605_1;
wire na606_1;
wire na607_1;
wire na608_1;
wire na609_1;
wire na610_1;
wire na611_1;
wire na612_1;
wire na613_1;
wire na614_1;
wire na615_1;
wire na616_1;
wire na617_1;
wire na618_1;
wire na619_1;
wire na620_1;
wire na621_1;
wire na622_1;
wire na623_1;
wire na624_1;
wire na625_1;
wire na626_1;
wire na627_1;
wire na628_1;
wire na629_1;
wire na630_1;
wire na631_1;
wire na632_1;
wire na633_1;
wire na634_1;
wire na635_1;
wire na636_1;
wire na637_1;
wire na638_1;
wire na639_1;
wire na640_1;
wire na641_1;
wire na642_1;
wire na643_1;
wire na644_1;
wire na645_1;
wire na646_1;
wire na647_1;
wire na648_1;
wire na649_1;
wire na650_1;
wire na651_1;
wire na652_1;
wire na653_1;
wire na654_1;
wire na655_1;
wire na656_1;
wire na657_1;
wire na658_1;
wire na659_1;
wire na660_1;
wire na661_1;
wire na662_1;
wire na663_1;
wire na664_1;
wire na665_1;
wire na666_1;
wire na667_1;
wire na668_1;
wire na669_1;
wire na670_1;
wire na671_1;
wire na672_1;
wire na673_1;
wire na674_1;
wire na675_1;
wire na676_1;
wire na677_1;
wire na678_1;
wire na679_1;
wire na680_1;
wire na681_1;
wire na682_1;
wire na683_1;
wire na684_1;
wire na685_1;
wire na686_1;
wire na687_1;
wire na688_1;
wire na689_1;
wire na690_1;
wire na691_1;
wire na692_1;
wire na693_1;
wire na694_1;
wire na695_1;
wire na696_1;
wire na697_1;
wire na698_1;
wire na699_1;
wire na700_1;
wire na701_1;
wire na702_1;
wire na703_1;
wire na704_1;
wire na705_1;
wire na706_1;
wire na707_1;
wire na708_1;
wire na709_1;
wire na710_1;
wire na711_1;
wire na712_1;
wire na713_1;
wire na714_1;
wire na715_1;
wire na716_1;
wire na717_1;
wire na718_1;
wire na719_1;
wire na720_1;
wire na721_1;
wire na722_1;
wire na723_1;
wire na724_1;
wire na725_1;
wire na726_1;
wire na727_1;
wire na728_1;
wire na729_1;
wire na730_1;
wire na731_1;
wire na732_1;
wire na733_1;
wire na734_1;
wire na735_1;
wire na736_1;
wire na737_1;
wire na738_1;
wire na739_1;
wire na740_1;
wire na741_1;
wire na742_1;
wire na743_1;
wire na744_1;
wire na745_1;
wire na746_1;
wire na747_1;
wire na748_1;
wire na749_1;
wire na750_1;
wire na751_1;
wire na752_1;
wire na753_1;
wire na754_1;
wire na755_1;
wire na756_1;
wire na757_1;
wire na758_1;
wire na759_1;
wire na760_1;
wire na761_1;
wire na762_1;
wire na763_1;
wire na764_1;
wire na765_1;
wire na766_1;
wire na767_1;
wire na768_1;
wire na769_1;
wire na770_1;
wire na771_1;
wire na772_1;
wire na773_1;
wire na774_1;
wire na775_1;
wire na776_1;
wire na777_1;
wire na778_1;
wire na779_1;
wire na780_1;
wire na781_1;
wire na782_1;
wire na783_1;
wire na784_1;
wire na785_1;
wire na786_1;
wire na787_1;
wire na788_1;
wire na789_1;
wire na790_1;
wire na791_1;
wire na792_1;
wire na793_1;
wire na794_1;
wire na795_1;
wire na796_1;
wire na797_1;
wire na798_1;
wire na799_1;
wire na800_2;
wire na801_1;
wire na802_2;
wire na803_1;
wire na804_2;
wire na805_1;
wire na806_2;
wire na807_1;
wire na808_2;
wire na809_1;
wire na810_1;
wire na811_1;
wire na812_2;
wire na813_1;
wire na814_1;
wire na815_2;
wire na816_2;
wire na817_1;
wire na818_1;
wire na819_1;
wire na822_1;
wire na823_1;
wire na824_1;
wire na826_2;
wire na827_1;
wire na828_2;
wire na829_1;
wire na830_1;
wire na831_1;
wire na832_1;
wire na833_1;
wire na834_1;
wire na835_1;
wire na836_2;
wire na837_1;
wire na838_1;
wire na840_1;
wire na841_1;
wire na842_2;
wire na843_1;
wire na844_1;
wire na845_2;
wire na846_1;
wire na847_1;
wire na848_1;
wire na849_1;
wire na850_1;
wire na851_1;
wire na852_1;
wire na853_1;
wire na854_1;
wire na855_1;
wire na856_2;
wire na857_1;
wire na858_1;
wire na859_2;
wire na861_1;
wire na862_2;
wire na863_2;
wire na864_1;
wire na865_1;
wire na866_2;
wire na867_1;
wire na868_2;
wire na869_1;
wire na870_1;
wire na871_1;
wire na872_1;
wire na873_1;
wire na874_1;
wire na875_2;
wire na876_1;
wire na877_2;
wire na878_1;
wire na879_2;
wire na880_1;
wire na881_1;
wire na883_1;
wire na884_1;
wire na885_2;
wire na886_1;
wire na887_1;
wire na888_1;
wire na889_1;
wire na890_2;
wire na891_1;
wire na892_2;
wire na893_2;
wire na894_2;
wire na896_1;
wire na897_1;
wire na899_1;
wire na900_1;
wire na901_1;
wire na902_1;
wire na903_1;
wire na904_1;
wire na905_1;
wire na906_1;
wire na907_1;
wire na908_1;
wire na909_2;
wire na911_2;
wire na912_1;
wire na913_1;
wire na914_1;
wire na915_1;
wire na916_1;
wire na917_1;
wire na918_2;
wire na919_2;
wire na920_1;
wire na921_1;
wire na922_1;
wire na923_1;
wire na924_1;
wire na925_1;
wire na926_1;
wire na928_1;
wire na929_1;
wire na930_1;
wire na931_1;
wire na932_1;
wire na933_1;
wire na934_1;
wire na935_1;
wire na936_1;
wire na937_2;
wire na938_1;
wire na939_2;
wire na940_1;
wire na941_1;
wire na942_2;
wire na943_2;
wire na944_2;
wire na945_1;
wire na946_1;
wire na947_1;
wire na948_2;
wire na949_2;
wire na951_1;
wire na952_2;
wire na953_1;
wire na954_1;
wire na955_1;
wire na956_1;
wire na957_2;
wire na958_1;
wire na959_1;
wire na961_1;
wire na962_1;
wire na963_2;
wire na964_1;
wire na965_2;
wire na966_2;
wire na967_1;
wire na968_1;
wire na969_1;
wire na970_1;
wire na973_1;
wire na974_1;
wire na975_1;
wire na977_1;
wire na978_2;
wire na979_1;
wire na980_1;
wire na981_1;
wire na982_1;
wire na983_1;
wire na984_1;
wire na985_1;
wire na986_2;
wire na987_1;
wire na988_1;
wire na989_2;
wire na990_1;
wire na991_1;
wire na992_2;
wire na993_1;
wire na994_1;
wire na995_2;
wire na996_2;
wire na997_1;
wire na998_1;
wire na999_1;
wire reset_n;
wire data_out;
wire na1000_1;
wire na1001_2;
wire na1002_1;
wire na1003_1;
wire na1005_1;
wire na1006_1;
wire na1007_1;
wire na1008_2;
wire na1009_1;
wire na1010_1;
wire na1011_1;
wire na1012_1;
wire na1013_2;
wire na1014_2;
wire na1015_1;
wire na1016_1;
wire na1018_1;
wire na1019_2;
wire na1020_1;
wire na1021_1;
wire na1022_1;
wire na1023_1;
wire na1024_1;
wire na1025_1;
wire na1026_2;
wire na1028_1;
wire na1029_1;
wire na1030_1;
wire na1031_1;
wire na1032_1;
wire na1033_1;
wire na1034_2;
wire na1035_1;
wire na1036_1;
wire na1037_1;
wire na1038_1;
wire na1039_1;
wire na1040_1;
wire na1041_1;
wire na1042_1;
wire na1043_1;
wire na1044_1;
wire na1045_1;
wire na1046_1;
wire na1047_1;
wire na1048_1;
wire na1049_1;
wire na1050_1;
wire na1051_1;
wire na1052_1;
wire na1053_1;
wire na1054_1;
wire na1055_1;
wire na1056_1;
wire na1057_1;
wire na1058_1;
wire na1059_1;
wire na1060_1;
wire na1061_1;
wire na1062_1;
wire na1063_1;
wire na1064_1;
wire na1065_1;
wire na1066_1;
wire na1067_1;
wire na1068_1;
wire na1069_1;
wire na1070_1;
wire na1071_1;
wire na1072_1;
wire na1073_1;
wire na1074_1;
wire na1075_1;
wire na1076_1;
wire na1077_1;
wire na1078_1;
wire na1079_1;
wire na1080_1;
wire na1081_1;
wire na1082_1;
wire na1083_1;
wire na1084_1;
wire na1085_1;
wire na1086_1;
wire na1087_1;
wire na1088_1;
wire na1089_1;
wire na1090_1;
wire na1091_1;
wire na1092_1;
wire na1093_1;
wire na1094_1;
wire na1095_1;
wire na1096_1;
wire na1097_1;
wire na1098_1;
wire na1099_1;
wire na1100_1;
wire na1101_1;
wire na1102_1;
wire na1103_1;
wire na1104_1;
wire na1105_1;
wire na1106_1;
wire na1107_1;
wire na1108_1;
wire na1109_1;
wire na1110_1;
wire na1111_1;
wire na1112_1;
wire na1113_1;
wire na1114_1;
wire na1115_1;
wire na1116_1;
wire na1117_1;
wire na1118_1;
wire na1119_1;
wire na1120_1;
wire na1121_1;
wire na1122_1;
wire na1123_1;
wire na1124_1;
wire na1125_1;
wire na1126_2;
wire na1127_1;
wire na1128_1;
wire na1129_1;
wire na1130_1;
wire na1131_1;
wire na1132_1;
wire na1133_1;
wire na1134_1;
wire na1135_1;
wire na1136_2;
wire na1137_1;
wire na1138_1;
wire na1139_1;
wire na1140_1;
wire na1141_1;
wire na1142_1;
wire na1143_1;
wire na1144_1;
wire na1145_1;
wire na1146_1;
wire na1147_1;
wire na1148_1;
wire na1149_1;
wire na1150_1;
wire na1151_1;
wire na1152_1;
wire na1153_1;
wire na1154_1;
wire na1155_1;
wire na1156_1;
wire na1157_1;
wire na1158_1;
wire na1159_1;
wire na1160_1;
wire na1161_1;
wire na1162_1;
wire na1163_1;
wire na1164_1;
wire na1165_1;
wire na1166_1;
wire na1167_1;
wire na1168_1;
wire na1169_1;
wire na1170_1;
wire na1171_1;
wire na1172_1;
wire na1173_1;
wire na1174_1;
wire na1175_1;
wire na1176_1;
wire na1177_1;
wire na1178_1;
wire na1179_1;
wire na1180_1;
wire na1181_1;
wire na1182_1;
wire na1183_1;
wire na1184_1;
wire na1185_1;
wire na1186_1;
wire na1187_1;
wire na1188_1;
wire na1189_1;
wire na1190_1;
wire na1191_1;
wire na1192_1;
wire na1193_1;
wire na1194_1;
wire na1195_1;
wire na1196_1;
wire na1197_1;
wire na1198_1;
wire na1199_1;
wire na1200_1;
wire na1201_2;
wire na1202_1;
wire na1203_1;
wire na1206_2;
wire na1207_2;
wire na1208_1;
wire na1209_1;
wire na1211_2;
wire na1212_1;
wire na1213_2;
wire na1214_1;
wire na1217_1;
wire na1219_2;
wire na1220_1;
wire na1222_2;
wire na1223_1;
wire na1224_2;
wire na1226_2;
wire na1227_1;
wire na1229_2;
wire na1230_2;
wire na1232_1;
wire na1233_2;
wire na1235_1;
wire na1236_2;
wire na1237_1;
wire na1239_1;
wire na1242_2;
wire na1243_1;
wire na1244_1;
wire na1245_2;
wire na1248_1;
wire na1251_2;
wire na1254_1;
wire na1255_1;
wire na1260_1;
wire na1262_2;
wire na1265_2;
wire na1266_1;
wire na1267_1;
wire na1268_2;
wire na1271_1;
wire na1276_1;
wire na1277_1;
wire na1282_1;
wire na1287_1;
wire na1288_1;
wire na1293_1;
wire na1295_1;
wire na1298_2;
wire na1299_1;
wire na1300_2;
wire na1301_2;
wire na1304_1;
wire na1306_2;
wire na1309_1;
wire na1312_2;
wire na1313_1;
wire na1316_1;
wire na1317_1;
wire na1318_1;
wire na1319_1;
wire na1320_2;
wire na1321_1;
wire na1322_2;
wire na1323_1;
wire na1324_2;
wire na1325_1;
wire na1328_2;
wire na1329_1;
wire na1330_2;
wire na1331_1;
wire na1332_2;
wire na1333_1;
wire na1334_1;
wire na1336_2;
wire na1337_1;
wire na1338_2;
wire na1339_1;
wire na1340_1;
wire na1341_1;
wire na1342_2;
wire na1343_1;
wire na1344_2;
wire na1345_1;
wire na1346_2;
wire na1347_1;
wire na1348_1;
wire na1349_1;
wire na1350_1;
wire na1351_1;
wire na1352_1;
wire na1353_1;
wire na1354_1;
wire na1355_1;
wire na1356_2;
wire na1357_1;
wire na1358_1;
wire na1361_1;
wire na1362_1;
wire na1363_2;
wire na1364_1;
wire na1365_2;
wire na1366_1;
wire na1367_2;
wire na1368_1;
wire na1369_2;
wire na1370_1;
wire na1371_2;
wire na1372_1;
wire na1373_2;
wire na1374_1;
wire na1375_1;
wire na1376_1;
wire na1377_2;
wire na1378_1;
wire na1379_2;
wire na1380_1;
wire na1381_1;
wire na1382_2;
wire na1383_1;
wire na1384_1;
wire na1385_1;
wire na1386_2;
wire na1387_1;
wire na1388_2;
wire na1389_1;
wire na1390_2;
wire na1391_1;
wire na1392_2;
wire na1393_2;
wire na1394_1;
wire na1395_1;
wire na1396_1;
wire na1397_2;
wire na1398_2;
wire na1399_1;
wire na1400_2;
wire na1401_2;
wire na1402_1;
wire na1403_2;
wire na1404_1;
wire na1405_2;
wire na1406_1;
wire na1407_2;
wire na1408_2;
wire na1409_1;
wire na1410_2;
wire na1411_1;
wire na1412_2;
wire na1413_2;
wire na1414_1;
wire na1415_1;
wire na1416_2;
wire na1417_1;
wire na1418_2;
wire na1419_2;
wire na1420_1;
wire na1421_1;
wire na1422_2;
wire na1423_2;
wire na1424_2;
wire na1425_2;
wire na1426_1;
wire na1427_2;
wire na1428_2;
wire na1429_1;
wire na1430_1;
wire na1431_2;
wire na1432_1;
wire na1433_2;
wire na1434_1;
wire na1435_2;
wire na1436_1;
wire na1437_2;
wire na1438_2;
wire na1439_2;
wire na1440_1;
wire na1441_2;
wire na1442_2;
wire na1443_1;
wire na1445_1;
wire na1446_1;
wire na1447_2;
wire na1449_1;
wire na1450_1;
wire na1451_1;
wire na1452_1;
wire na1453_1;
wire na1454_1;
wire na1455_2;
wire na1456_1;
wire na1457_1;
wire na1458_2;
wire na1459_1;
wire na1460_1;
wire na1461_2;
wire na1462_1;
wire na1464_2;
wire na1465_1;
wire na1466_2;
wire na1467_2;
wire na1468_1;
wire na1469_1;
wire na1470_1;
wire na1471_1;
wire na1473_1;
wire na1475_2;
wire na1476_1;
wire na1477_1;
wire na1478_1;
wire na1480_1;
wire na1481_2;
wire na1482_1;
wire na1483_2;
wire na1484_1;
wire na1485_1;
wire na1486_1;
wire na1487_2;
wire na1488_2;
wire na1489_2;
wire na1490_2;
wire na1491_2;
wire na1492_1;
wire na1493_2;
wire na1494_1;
wire na1495_2;
wire na1496_1;
wire na1497_2;
wire na1498_2;
wire na1499_1;
wire na1500_1;
wire na1501_2;
wire na1502_1;
wire na1503_1;
wire na1504_1;
wire na1505_2;
wire na1506_1;
wire na1507_2;
wire na1508_1;
wire na1509_2;
wire na1510_1;
wire na1511_2;
wire na1512_2;
wire na1513_1;
wire na1514_2;
wire na1515_1;
wire na1516_2;
wire na1517_2;
wire na1518_2;
wire na1519_1;
wire na1520_1;
wire na1521_2;
wire na1522_1;
wire na1523_1;
wire na1524_2;
wire na1525_1;
wire na1526_1;
wire na1527_1;
wire na1528_2;
wire na1529_2;
wire na1530_2;
wire na1531_2;
wire na1532_2;
wire na1533_1;
wire na1534_1;
wire na1535_1;
wire na1536_2;
wire na1537_1;
wire na1538_2;
wire na1539_1;
wire na1540_2;
wire na1541_1;
wire na1542_1;
wire na1543_1;
wire na1544_2;
wire na1545_1;
wire na1546_2;
wire na1547_1;
wire na1548_1;
wire na1549_1;
wire na1550_1;
wire na1551_2;
wire na1552_1;
wire na1553_2;
wire na1554_1;
wire na1555_2;
wire na1556_2;
wire na1557_1;
wire na1558_2;
wire na1559_1;
wire na1560_2;
wire na1561_1;
wire na1562_1;
wire na1563_2;
wire na1564_1;
wire na1565_2;
wire na1566_2;
wire na1567_1;
wire na1568_2;
wire na1569_2;
wire na1570_1;
wire na1571_2;
wire na1572_1;
wire na1573_2;
wire na1574_1;
wire na1575_1;
wire na1576_2;
wire na1577_1;
wire na1578_1;
wire na1579_1;
wire na1580_1;
wire na1581_1;
wire na1582_1;
wire na1583_2;
wire na1584_1;
wire na1585_1;
wire na1586_1;
wire na1587_2;
wire na1588_2;
wire na1589_1;
wire na1590_1;
wire na1591_2;
wire na1592_1;
wire na1593_2;
wire na1594_1;
wire na1595_2;
wire na1596_1;
wire na1597_2;
wire na1598_1;
wire na1599_1;
wire na1600_1;
wire na1601_2;
wire na1602_1;
wire na1603_2;
wire na1604_2;
wire na1605_2;
wire na1606_1;
wire na1607_2;
wire na1608_2;
wire na1609_2;
wire na1610_1;
wire na1611_2;
wire na1612_1;
wire na1613_1;
wire na1614_2;
wire na1615_2;
wire na1616_1;
wire na1617_2;
wire na1618_1;
wire na1619_1;
wire na1620_1;
wire na1621_2;
wire na1622_2;
wire na1623_1;
wire na1624_1;
wire na1625_2;
wire na1626_1;
wire na1627_2;
wire na1628_2;
wire na1629_2;
wire na1630_1;
wire na1631_2;
wire na1632_1;
wire na1633_1;
wire na1634_2;
wire na1635_2;
wire na1636_1;
wire na1637_1;
wire na1638_2;
wire na1639_1;
wire na1640_2;
wire na1641_2;
wire na1642_1;
wire na1643_1;
wire na1644_1;
wire na1645_1;
wire na1646_1;
wire na1647_2;
wire na1648_2;
wire na1649_2;
wire na1650_1;
wire na1651_2;
wire na1652_1;
wire na1653_2;
wire na1654_2;
wire na1655_2;
wire na1656_1;
wire na1657_1;
wire na1658_2;
wire na1659_2;
wire na1660_1;
wire na1661_2;
wire na1662_2;
wire na1663_2;
wire na1664_1;
wire na1665_2;
wire na1666_1;
wire na1667_2;
wire na1668_1;
wire na1669_2;
wire na1670_2;
wire na1671_2;
wire na1672_2;
wire na1673_2;
wire na1674_1;
wire na1675_2;
wire na1676_2;
wire na1677_2;
wire na1678_2;
wire na1679_1;
wire na1680_1;
wire na1681_2;
wire na1682_2;
wire na1683_1;
wire na1684_1;
wire na1685_1;
wire na1686_1;
wire na1687_2;
wire na1688_1;
wire na1689_2;
wire na1690_2;
wire na1691_1;
wire na1692_1;
wire na1693_2;
wire na1694_2;
wire na1695_1;
wire na1696_1;
wire na1697_2;
wire na1698_1;
wire na1699_2;
wire na1700_1;
wire na1701_2;
wire na1702_1;
wire na1703_1;
wire na1704_1;
wire na1705_1;
wire na1706_2;
wire na1707_2;
wire na1708_1;
wire na1709_1;
wire na1710_2;
wire na1711_1;
wire na1712_1;
wire na1713_1;
wire na1714_2;
wire na1715_1;
wire na1716_2;
wire na1717_1;
wire na1718_1;
wire na1719_1;
wire na1720_2;
wire na1721_1;
wire na1722_1;
wire na1723_1;
wire na1724_2;
wire na1725_2;
wire na1726_1;
wire na1727_1;
wire na1728_1;
wire na1729_1;
wire na1730_1;
wire na1731_1;
wire na1732_2;
wire na1733_1;
wire na1735_1;
wire na1737_1;
wire na1739_1;
wire na1741_1;
wire na1743_1;
wire na1745_2;
wire na1746_1;
wire na1747_1;
wire na1748_1;
wire na1750_1;
wire na1752_1;
wire na1754_1;
wire na1756_1;
wire na1758_1;
wire na1760_2;
wire na1761_1;
wire na1763_1;
wire na1765_1;
wire na1767_1;
wire na1769_1;
wire na1770_1;
wire na1771_1;
wire na1773_1;
wire na1775_1;
wire na1776_2;
wire na1777_1;
wire na1779_1;
wire na1781_1;
wire na1783_1;
wire na1784_1;
wire na1797_1;
wire na1799_1;
wire na1800_1;
wire na1801_1;
wire na1803_1;
wire na1804_2;
wire na1805_1;
wire na1806_1;
wire na1808_1;
wire na1809_1;
wire na1810_1;
wire na1811_1;
wire na1813_1;
wire na1814_2;
wire na1815_1;
wire na1816_1;
wire na1818_1;
wire na1819_1;
wire na1820_1;
wire na1821_1;
wire na1823_1;
wire na1824_2;
wire na1825_1;
wire na1826_1;
wire na1828_1;
wire na1829_2;
wire na1830_1;
wire na1831_1;
wire na1832_1;
wire na1833_2;
wire na1834_1;
wire na1835_1;
wire na1836_2;
wire na1837_1;
wire na1838_1;
wire na1839_1;
wire na1840_1;
wire na1841_1;
wire na1842_1;
wire na1843_2;
wire na1844_2;
wire na1845_1;
wire na1846_2;
wire na1847_1;
wire na1848_1;
wire na1849_1;
wire na1850_1;
wire na1852_4;
wire na1854_4;
wire na1856_4;
wire na1858_4;
wire na1859_1;
wire na1859_4;
wire na1860_1;
wire na1860_2;
wire na1860_4;
wire na1862_1;
wire na1862_2;
wire na1862_4;
wire na1864_1;
wire na1865_1;
wire na1865_4;
wire na1866_1;
wire na1866_2;
wire na1866_4;
wire na1868_1;
wire na1868_2;
wire na1870_1;
wire na1870_4;
wire na1871_1;
wire na1871_2;
wire na1871_4;
wire na1873_1;
wire na1874_1;
wire na1874_4;
wire na1876_1;
wire na1876_2;
wire na1876_4;
wire na1878_1;
wire na1878_2;
wire na1878_4;
wire na1880_1;
wire na1880_2;
wire na1880_4;
wire na1882_1;
wire na1882_2;
wire na1882_4;
wire na1884_1;
wire na1884_2;
wire na1885_1;
wire na1885_4;
wire na1886_1;
wire na1886_2;
wire na1888_1;
wire na1888_4;
wire na1890_1;
wire na1890_2;
wire na1890_4;
wire na1892_1;
wire na1892_2;
wire na1892_4;
wire na1894_1;
wire na1894_2;
wire na1894_4;
wire na1896_1;
wire na1896_2;
wire na1896_4;
wire na1898_1;
wire na1898_2;
wire na1899_1;
wire na1899_4;
wire na1900_1;
wire na1900_2;
wire na1903_2;
wire na1903_2_i;
wire na1904_1;
wire na1904_1_i;
wire na1905_2;
wire na1905_2_i;
wire na1906_1;
wire na1906_1_i;
wire na1907_2;
wire na1907_2_i;
wire na1908_1;
wire na1908_1_i;
wire na1909_2;
wire na1909_2_i;
wire na1910_1;
wire na1910_1_i;
wire na1911_2;
wire na1911_2_i;
wire na1912_1;
wire na1912_1_i;
wire na1913_2;
wire na1913_2_i;
wire na1914_1;
wire na1914_1_i;
wire na1915_2;
wire na1915_2_i;
wire na1916_1;
wire na1916_1_i;
wire na1917_2;
wire na1917_2_i;
wire na1918_1;
wire na1918_1_i;
wire na1919_2;
wire na1919_2_i;
wire na1920_1;
wire na1920_1_i;
wire na1921_2;
wire na1921_2_i;
wire na1922_1;
wire na1922_1_i;
wire na1923_2;
wire na1923_2_i;
wire na1924_1;
wire na1924_1_i;
wire na1925_2;
wire na1925_2_i;
wire na1926_1;
wire na1926_1_i;
wire na1927_2;
wire na1927_2_i;
wire na1928_1;
wire na1929_1;
wire na1929_1_i;
wire na1930_1;
wire na1930_1_i;
wire na1930_2;
wire na1930_2_i;
wire na1932_1;
wire na1932_1_i;
wire na1932_2;
wire na1932_2_i;
wire na1934_2;
wire na1934_2_i;
wire na1935_1;
wire na1935_1_i;
wire na1935_2;
wire na1935_2_i;
wire na1937_1;
wire na1937_1_i;
wire na1937_2;
wire na1937_2_i;
wire na1938_1;
wire na1938_1_i;
wire na1941_1;
wire na1941_1_i;
wire na1941_2;
wire na1941_2_i;
wire na1943_1;
wire na1943_1_i;
wire na1943_2;
wire na1943_2_i;
wire na1945_1;
wire na1945_1_i;
wire na1945_2;
wire na1945_2_i;
wire na1946_1;
wire na1946_1_i;
wire na1946_2;
wire na1946_2_i;
wire na1947_2;
wire na1947_2_i;
wire na1948_1;
wire na1948_1_i;
wire na1949_2;
wire na1949_2_i;
wire na1950_1;
wire na1950_1_i;
wire na1951_2;
wire na1951_2_i;
wire na1952_1;
wire na1952_1_i;
wire na1953_2;
wire na1953_2_i;
wire na1954_1;
wire na1954_1_i;
wire na1955_2;
wire na1955_2_i;
wire na1956_1;
wire na1956_1_i;
wire na1957_2;
wire na1957_2_i;
wire na1958_1;
wire na1958_1_i;
wire na1959_2;
wire na1959_2_i;
wire na1960_1;
wire na1960_1_i;
wire na1961_2;
wire na1961_2_i;
wire na1962_1;
wire na1962_1_i;
wire na1963_2;
wire na1963_2_i;
wire na1964_1;
wire na1964_1_i;
wire na1965_2;
wire na1965_2_i;
wire na1966_1;
wire na1966_1_i;
wire na1967_2;
wire na1967_2_i;
wire na1968_1;
wire na1968_1_i;
wire na1969_2;
wire na1969_2_i;
wire na1970_1;
wire na1970_1_i;
wire na1971_2;
wire na1971_2_i;
wire na1972_1;
wire na1972_1_i;
wire na1973_2;
wire na1973_2_i;
wire na1974_1;
wire na1974_1_i;
wire na1975_2;
wire na1975_2_i;
wire na1976_1;
wire na1976_1_i;
wire na1977_2;
wire na1977_2_i;
wire na1978_1;
wire na1978_1_i;
wire na1979_2;
wire na1979_2_i;
wire na1980_1;
wire na1980_1_i;
wire na1981_2;
wire na1981_2_i;
wire na1982_1;
wire na1982_1_i;
wire na1983_2;
wire na1983_2_i;
wire na1984_1;
wire na1984_1_i;
wire na1985_2;
wire na1985_2_i;
wire na1986_1;
wire na1986_1_i;
wire na1987_2;
wire na1987_2_i;
wire na1988_1;
wire na1988_1_i;
wire na1989_2;
wire na1989_2_i;
wire na1990_1;
wire na1990_1_i;
wire na1991_1;
wire na1991_1_i;
wire na1992_1;
wire na1992_1_i;
wire na1993_2;
wire na1993_2_i;
wire na1994_1;
wire na1994_1_i;
wire na1995_2;
wire na1995_2_i;
wire na1996_1;
wire na1996_1_i;
wire na1997_2;
wire na1997_2_i;
wire na1998_1;
wire na1998_1_i;
wire na1999_2;
wire na1999_2_i;
wire na2000_1;
wire na2000_1_i;
wire na2001_2;
wire na2001_2_i;
wire na2002_1;
wire na2002_1_i;
wire na2003_2;
wire na2003_2_i;
wire na2004_1;
wire na2004_1_i;
wire na2005_2;
wire na2005_2_i;
wire na2006_1;
wire na2006_1_i;
wire na2007_2;
wire na2007_2_i;
wire na2008_1;
wire na2008_1_i;
wire na2009_2;
wire na2009_2_i;
wire na2010_1;
wire na2010_1_i;
wire na2011_2;
wire na2011_2_i;
wire na2012_1;
wire na2012_1_i;
wire na2013_2;
wire na2013_2_i;
wire na2014_1;
wire na2014_1_i;
wire na2015_2;
wire na2015_2_i;
wire na2016_1;
wire na2016_1_i;
wire na2017_2;
wire na2017_2_i;
wire na2018_1;
wire na2018_1_i;
wire na2019_2;
wire na2019_2_i;
wire na2020_1;
wire na2020_1_i;
wire na2021_2;
wire na2021_2_i;
wire na2022_1;
wire na2022_1_i;
wire na2023_2;
wire na2023_2_i;
wire na2024_1;
wire na2024_1_i;
wire na2025_2;
wire na2025_2_i;
wire na2026_1;
wire na2026_1_i;
wire na2027_2;
wire na2027_2_i;
wire na2028_1;
wire na2028_1_i;
wire na2029_2;
wire na2029_2_i;
wire na2030_1;
wire na2030_1_i;
wire na2031_2;
wire na2031_2_i;
wire na2032_1;
wire na2032_1_i;
wire na2033_2;
wire na2033_2_i;
wire na2034_1;
wire na2034_1_i;
wire na2035_2;
wire na2035_2_i;
wire na2036_1;
wire na2036_1_i;
wire na2037_2;
wire na2037_2_i;
wire na2038_1;
wire na2038_1_i;
wire na2039_2;
wire na2039_2_i;
wire na2040_1;
wire na2040_1_i;
wire na2041_2;
wire na2041_2_i;
wire na2042_1;
wire na2042_1_i;
wire na2043_2;
wire na2043_2_i;
wire na2044_1;
wire na2044_1_i;
wire na2045_2;
wire na2045_2_i;
wire na2046_1;
wire na2046_1_i;
wire na2047_2;
wire na2047_2_i;
wire na2048_1;
wire na2048_1_i;
wire na2049_2;
wire na2049_2_i;
wire na2050_1;
wire na2050_1_i;
wire na2051_2;
wire na2051_2_i;
wire na2052_1;
wire na2052_1_i;
wire na2053_2;
wire na2053_2_i;
wire na2054_1;
wire na2054_1_i;
wire na2055_2;
wire na2055_2_i;
wire na2056_1;
wire na2056_1_i;
wire na2057_2;
wire na2057_2_i;
wire na2058_1;
wire na2058_1_i;
wire na2059_2;
wire na2059_2_i;
wire na2060_1;
wire na2060_1_i;
wire na2061_2;
wire na2061_2_i;
wire na2062_1;
wire na2062_1_i;
wire na2063_2;
wire na2063_2_i;
wire na2064_1;
wire na2064_1_i;
wire na2065_2;
wire na2065_2_i;
wire na2066_1;
wire na2066_1_i;
wire na2067_2;
wire na2067_2_i;
wire na2068_1;
wire na2068_1_i;
wire na2069_2;
wire na2069_2_i;
wire na2070_1;
wire na2070_1_i;
wire na2071_2;
wire na2071_2_i;
wire na2072_1;
wire na2072_1_i;
wire na2073_2;
wire na2073_2_i;
wire na2074_1;
wire na2074_1_i;
wire na2075_2;
wire na2075_2_i;
wire na2076_1;
wire na2076_1_i;
wire na2077_2;
wire na2077_2_i;
wire na2078_1;
wire na2078_1_i;
wire na2079_2;
wire na2079_2_i;
wire na2080_1;
wire na2080_1_i;
wire na2081_2;
wire na2081_2_i;
wire na2082_1;
wire na2082_1_i;
wire na2083_2;
wire na2083_2_i;
wire na2084_1;
wire na2084_1_i;
wire na2085_2;
wire na2085_2_i;
wire na2086_1;
wire na2086_1_i;
wire na2087_2;
wire na2087_2_i;
wire na2088_1;
wire na2088_1_i;
wire na2089_2;
wire na2089_2_i;
wire na2090_1;
wire na2090_1_i;
wire na2091_2;
wire na2091_2_i;
wire na2092_1;
wire na2092_1_i;
wire na2093_2;
wire na2093_2_i;
wire na2094_1;
wire na2094_1_i;
wire na2095_2;
wire na2095_2_i;
wire na2096_1;
wire na2096_1_i;
wire na2097_2;
wire na2097_2_i;
wire na2098_1;
wire na2098_1_i;
wire na2099_2;
wire na2099_2_i;
wire na2100_1;
wire na2100_1_i;
wire na2101_2;
wire na2101_2_i;
wire na2102_1;
wire na2102_1_i;
wire na2103_2;
wire na2103_2_i;
wire na2104_1;
wire na2104_1_i;
wire na2105_2;
wire na2105_2_i;
wire na2106_1;
wire na2106_1_i;
wire na2107_2;
wire na2107_2_i;
wire na2108_1;
wire na2108_1_i;
wire na2109_2;
wire na2109_2_i;
wire na2110_1;
wire na2110_1_i;
wire na2111_2;
wire na2111_2_i;
wire na2112_1;
wire na2112_1_i;
wire na2113_2;
wire na2113_2_i;
wire na2114_1;
wire na2114_1_i;
wire na2115_2;
wire na2115_2_i;
wire na2116_1;
wire na2116_1_i;
wire na2117_2;
wire na2117_2_i;
wire na2118_1;
wire na2118_1_i;
wire na2119_2;
wire na2119_2_i;
wire na2120_1;
wire na2120_1_i;
wire na2121_2;
wire na2121_2_i;
wire na2122_1;
wire na2122_1_i;
wire na2123_2;
wire na2123_2_i;
wire na2124_1;
wire na2124_1_i;
wire na2125_2;
wire na2125_2_i;
wire na2126_1;
wire na2126_1_i;
wire na2127_2;
wire na2127_2_i;
wire na2128_1;
wire na2128_1_i;
wire na2129_2;
wire na2129_2_i;
wire na2130_1;
wire na2130_1_i;
wire na2131_2;
wire na2131_2_i;
wire na2132_1;
wire na2132_1_i;
wire na2133_2;
wire na2133_2_i;
wire na2134_1;
wire na2134_1_i;
wire na2135_2;
wire na2135_2_i;
wire na2136_2;
wire na2136_2_i;
wire na2137_2;
wire na2137_2_i;
wire na2138_1;
wire na2138_1_i;
wire na2139_2;
wire na2139_2_i;
wire na2140_1;
wire na2140_1_i;
wire na2141_2;
wire na2141_2_i;
wire na2142_1;
wire na2142_1_i;
wire na2143_2;
wire na2143_2_i;
wire na2144_1;
wire na2144_1_i;
wire na2145_2;
wire na2145_2_i;
wire na2146_1;
wire na2146_1_i;
wire na2147_2;
wire na2147_2_i;
wire na2148_1;
wire na2148_1_i;
wire na2149_2;
wire na2149_2_i;
wire na2150_1;
wire na2150_1_i;
wire na2151_2;
wire na2151_2_i;
wire na2152_1;
wire na2152_1_i;
wire na2153_2;
wire na2153_2_i;
wire na2154_1;
wire na2154_1_i;
wire na2155_2;
wire na2155_2_i;
wire na2156_1;
wire na2156_1_i;
wire na2157_2;
wire na2157_2_i;
wire na2158_1;
wire na2158_1_i;
wire na2159_2;
wire na2159_2_i;
wire na2160_1;
wire na2160_1_i;
wire na2161_2;
wire na2161_2_i;
wire na2162_1;
wire na2162_1_i;
wire na2163_2;
wire na2163_2_i;
wire na2164_1;
wire na2164_1_i;
wire na2165_2;
wire na2165_2_i;
wire na2166_1;
wire na2166_1_i;
wire na2167_2;
wire na2167_2_i;
wire na2168_1;
wire na2168_1_i;
wire na2169_2;
wire na2169_2_i;
wire na2170_1;
wire na2170_1_i;
wire na2171_2;
wire na2171_2_i;
wire na2172_1;
wire na2172_1_i;
wire na2173_2;
wire na2173_2_i;
wire na2174_1;
wire na2174_1_i;
wire na2175_2;
wire na2175_2_i;
wire na2176_1;
wire na2176_1_i;
wire na2177_2;
wire na2177_2_i;
wire na2178_1;
wire na2178_1_i;
wire na2179_2;
wire na2179_2_i;
wire na2180_1;
wire na2180_1_i;
wire na2181_2;
wire na2181_2_i;
wire na2182_1;
wire na2182_1_i;
wire na2183_2;
wire na2183_2_i;
wire na2184_1;
wire na2184_1_i;
wire na2185_2;
wire na2185_2_i;
wire na2186_1;
wire na2186_1_i;
wire na2187_2;
wire na2187_2_i;
wire na2188_1;
wire na2188_1_i;
wire na2189_2;
wire na2189_2_i;
wire na2190_1;
wire na2190_1_i;
wire na2191_2;
wire na2191_2_i;
wire na2192_1;
wire na2192_1_i;
wire na2193_2;
wire na2193_2_i;
wire na2194_1;
wire na2194_1_i;
wire na2195_2;
wire na2195_2_i;
wire na2196_1;
wire na2196_1_i;
wire na2197_2;
wire na2197_2_i;
wire na2198_1;
wire na2198_1_i;
wire na2199_2;
wire na2199_2_i;
wire na2200_1;
wire na2200_1_i;
wire na2201_2;
wire na2201_2_i;
wire na2202_1;
wire na2202_1_i;
wire na2203_2;
wire na2203_2_i;
wire na2204_1;
wire na2204_1_i;
wire na2205_2;
wire na2205_2_i;
wire na2206_1;
wire na2206_1_i;
wire na2207_2;
wire na2207_2_i;
wire na2208_1;
wire na2208_1_i;
wire na2209_2;
wire na2209_2_i;
wire na2210_2;
wire na2210_2_i;
wire na2211_1;
wire na2211_1_i;
wire na2212_2;
wire na2212_2_i;
wire na2213_1;
wire na2213_1_i;
wire na2214_2;
wire na2214_2_i;
wire na2215_1;
wire na2215_1_i;
wire na2216_2;
wire na2216_2_i;
wire na2217_1;
wire na2217_1_i;
wire na2218_2;
wire na2218_2_i;
wire na2219_1;
wire na2219_1_i;
wire na2220_2;
wire na2220_2_i;
wire na2221_1;
wire na2221_1_i;
wire na2222_2;
wire na2222_2_i;
wire na2223_1;
wire na2223_1_i;
wire na2224_1;
wire na2224_1_i;
wire na2225_1;
wire na2225_1_i;
wire na2226_2;
wire na2226_2_i;
wire na2227_1;
wire na2227_1_i;
wire na2228_2;
wire na2228_2_i;
wire na2229_1;
wire na2229_1_i;
wire na2230_2;
wire na2230_2_i;
wire na2231_1;
wire na2231_1_i;
wire na2232_2;
wire na2232_2_i;
wire na2233_1;
wire na2233_1_i;
wire na2234_2;
wire na2234_2_i;
wire na2235_1;
wire na2235_1_i;
wire na2236_2;
wire na2236_2_i;
wire na2237_1;
wire na2237_1_i;
wire na2238_2;
wire na2238_2_i;
wire na2239_1;
wire na2239_1_i;
wire na2240_2;
wire na2240_2_i;
wire na2241_1;
wire na2241_1_i;
wire na2242_2;
wire na2242_2_i;
wire na2243_1;
wire na2243_1_i;
wire na2244_2;
wire na2244_2_i;
wire na2245_1;
wire na2245_1_i;
wire na2246_2;
wire na2246_2_i;
wire na2247_1;
wire na2247_1_i;
wire na2248_2;
wire na2248_2_i;
wire na2249_1;
wire na2249_1_i;
wire na2250_2;
wire na2250_2_i;
wire na2251_1;
wire na2251_1_i;
wire na2252_2;
wire na2252_2_i;
wire na2253_2;
wire na2253_2_i;
wire na2254_2;
wire na2254_2_i;
wire na2255_1;
wire na2255_1_i;
wire na2256_2;
wire na2256_2_i;
wire na2257_1;
wire na2257_1_i;
wire na2258_2;
wire na2258_2_i;
wire na2259_1;
wire na2259_1_i;
wire na2260_2;
wire na2260_2_i;
wire na2261_1;
wire na2261_1_i;
wire na2262_2;
wire na2262_2_i;
wire na2263_1;
wire na2263_1_i;
wire na2264_2;
wire na2264_2_i;
wire na2265_1;
wire na2265_1_i;
wire na2266_2;
wire na2266_2_i;
wire na2267_1;
wire na2267_1_i;
wire na2268_2;
wire na2268_2_i;
wire na2269_1;
wire na2269_1_i;
wire na2270_2;
wire na2270_2_i;
wire na2271_1;
wire na2271_1_i;
wire na2272_2;
wire na2272_2_i;
wire na2273_1;
wire na2273_1_i;
wire na2274_2;
wire na2274_2_i;
wire na2275_1;
wire na2275_1_i;
wire na2276_2;
wire na2276_2_i;
wire na2277_1;
wire na2277_1_i;
wire na2278_2;
wire na2278_2_i;
wire na2279_1;
wire na2279_1_i;
wire na2280_2;
wire na2280_2_i;
wire na2281_1;
wire na2281_1_i;
wire na2282_2;
wire na2282_2_i;
wire na2283_2;
wire na2283_2_i;
wire na2284_2;
wire na2284_2_i;
wire na2285_1;
wire na2285_1_i;
wire na2286_2;
wire na2286_2_i;
wire na2287_1;
wire na2287_1_i;
wire na2288_2;
wire na2288_2_i;
wire na2289_1;
wire na2289_1_i;
wire na2290_2;
wire na2290_2_i;
wire na2291_1;
wire na2291_1_i;
wire na2292_2;
wire na2292_2_i;
wire na2293_1;
wire na2293_1_i;
wire na2294_2;
wire na2294_2_i;
wire na2295_1;
wire na2295_1_i;
wire na2296_2;
wire na2296_2_i;
wire na2297_1;
wire na2297_1_i;
wire na2298_2;
wire na2298_2_i;
wire na2299_1;
wire na2299_1_i;
wire na2300_2;
wire na2300_2_i;
wire na2301_1;
wire na2301_1_i;
wire na2302_2;
wire na2302_2_i;
wire na2303_1;
wire na2303_1_i;
wire na2304_2;
wire na2304_2_i;
wire na2305_1;
wire na2305_1_i;
wire na2306_2;
wire na2306_2_i;
wire na2307_1;
wire na2307_1_i;
wire na2308_2;
wire na2308_2_i;
wire na2309_1;
wire na2309_1_i;
wire na2310_2;
wire na2310_2_i;
wire na2311_1;
wire na2311_1_i;
wire na2312_1;
wire na2312_1_i;
wire na2313_1;
wire na2313_1_i;
wire na2314_2;
wire na2314_2_i;
wire na2315_1;
wire na2315_1_i;
wire na2316_2;
wire na2316_2_i;
wire na2317_1;
wire na2317_1_i;
wire na2318_2;
wire na2318_2_i;
wire na2319_1;
wire na2319_1_i;
wire na2320_2;
wire na2320_2_i;
wire na2321_1;
wire na2321_1_i;
wire na2322_2;
wire na2322_2_i;
wire na2323_1;
wire na2323_1_i;
wire na2324_2;
wire na2324_2_i;
wire na2325_1;
wire na2325_1_i;
wire na2326_2;
wire na2326_2_i;
wire na2327_1;
wire na2327_1_i;
wire na2328_2;
wire na2328_2_i;
wire na2329_1;
wire na2329_1_i;
wire na2330_2;
wire na2330_2_i;
wire na2331_1;
wire na2331_1_i;
wire na2332_2;
wire na2332_2_i;
wire na2333_1;
wire na2333_1_i;
wire na2334_2;
wire na2334_2_i;
wire na2335_1;
wire na2335_1_i;
wire na2336_2;
wire na2336_2_i;
wire na2337_1;
wire na2337_1_i;
wire na2338_2;
wire na2338_2_i;
wire na2339_1;
wire na2339_1_i;
wire na2340_2;
wire na2340_2_i;
wire na2341_1;
wire na2341_1_i;
wire na2342_1;
wire na2342_1_i;
wire na2343_1;
wire na2343_1_i;
wire na2344_2;
wire na2344_2_i;
wire na2345_1;
wire na2345_1_i;
wire na2346_2;
wire na2346_2_i;
wire na2347_1;
wire na2347_1_i;
wire na2348_2;
wire na2348_2_i;
wire na2349_1;
wire na2349_1_i;
wire na2350_2;
wire na2350_2_i;
wire na2351_1;
wire na2351_1_i;
wire na2352_2;
wire na2352_2_i;
wire na2353_1;
wire na2353_1_i;
wire na2354_2;
wire na2354_2_i;
wire na2355_1;
wire na2355_1_i;
wire na2356_2;
wire na2356_2_i;
wire na2357_1;
wire na2357_1_i;
wire na2358_2;
wire na2358_2_i;
wire na2359_1;
wire na2359_1_i;
wire na2360_2;
wire na2360_2_i;
wire na2361_1;
wire na2361_1_i;
wire na2362_2;
wire na2362_2_i;
wire na2363_1;
wire na2363_1_i;
wire na2364_2;
wire na2364_2_i;
wire na2365_1;
wire na2365_1_i;
wire na2366_2;
wire na2366_2_i;
wire na2367_1;
wire na2367_1_i;
wire na2368_2;
wire na2368_2_i;
wire na2369_1;
wire na2369_1_i;
wire na2370_2;
wire na2370_2_i;
wire na2371_2;
wire na2371_2_i;
wire na2372_2;
wire na2372_2_i;
wire na2373_1;
wire na2373_1_i;
wire na2374_2;
wire na2374_2_i;
wire na2375_1;
wire na2375_1_i;
wire na2376_2;
wire na2376_2_i;
wire na2377_1;
wire na2377_1_i;
wire na2378_2;
wire na2378_2_i;
wire na2379_1;
wire na2379_1_i;
wire na2380_2;
wire na2380_2_i;
wire na2381_1;
wire na2381_1_i;
wire na2382_2;
wire na2382_2_i;
wire na2383_1;
wire na2383_1_i;
wire na2384_2;
wire na2384_2_i;
wire na2385_1;
wire na2385_1_i;
wire na2386_2;
wire na2386_2_i;
wire na2387_1;
wire na2387_1_i;
wire na2388_2;
wire na2388_2_i;
wire na2389_1;
wire na2389_1_i;
wire na2390_2;
wire na2390_2_i;
wire na2391_1;
wire na2391_1_i;
wire na2392_2;
wire na2392_2_i;
wire na2393_1;
wire na2393_1_i;
wire na2394_2;
wire na2394_2_i;
wire na2395_1;
wire na2395_1_i;
wire na2396_2;
wire na2396_2_i;
wire na2397_1;
wire na2397_1_i;
wire na2398_2;
wire na2398_2_i;
wire na2399_1;
wire na2399_1_i;
wire na2400_2;
wire na2400_2_i;
wire na2401_2;
wire na2401_2_i;
wire na2402_2;
wire na2402_2_i;
wire na2403_1;
wire na2403_1_i;
wire na2404_2;
wire na2404_2_i;
wire na2405_1;
wire na2405_1_i;
wire na2406_2;
wire na2406_2_i;
wire na2407_1;
wire na2407_1_i;
wire na2408_2;
wire na2408_2_i;
wire na2409_1;
wire na2409_1_i;
wire na2410_2;
wire na2410_2_i;
wire na2411_1;
wire na2411_1_i;
wire na2412_2;
wire na2412_2_i;
wire na2413_1;
wire na2413_1_i;
wire na2415_2;
wire na2415_2_i;
wire na2416_1;
wire na2416_1_i;
wire na2416_2;
wire na2416_2_i;
wire na2417_1;
wire na2417_1_i;
wire na2418_2;
wire na2418_2_i;
wire na2419_1;
wire na2419_1_i;
wire na2420_2;
wire na2420_2_i;
wire na2421_1;
wire na2421_1_i;
wire na2422_2;
wire na2422_2_i;
wire na2423_1;
wire na2423_1_i;
wire na2424_1;
wire na2424_1_i;
wire na2424_2;
wire na2424_2_i;
wire na2425_2;
wire na2425_2_i;
wire na2426_1;
wire na2426_1_i;
wire na2427_1;
wire na2427_1_i;
wire na2427_2;
wire na2427_2_i;
wire na2428_2;
wire na2428_2_i;
wire na2429_1;
wire na2429_1_i;
wire na2430_2;
wire na2430_2_i;
wire na2431_1;
wire na2431_1_i;
wire na2431_2;
wire na2431_2_i;
wire na2432_1;
wire na2432_1_i;
wire na2433_2;
wire na2433_2_i;
wire na2434_1;
wire na2434_1_i;
wire na2434_2;
wire na2434_2_i;
wire na2435_1;
wire na2435_1_i;
wire na2435_2;
wire na2435_2_i;
wire na2436_1;
wire na2436_1_i;
wire na2437_1;
wire na2437_1_i;
wire na2438_1;
wire na2438_1_i;
wire na2439_2;
wire na2439_2_i;
wire na2440_1;
wire na2440_1_i;
wire na2440_2;
wire na2440_2_i;
wire na2441_1;
wire na2441_1_i;
wire na2442_2;
wire na2442_2_i;
wire na2443_1;
wire na2443_1_i;
wire na2444_2;
wire na2444_2_i;
wire na2445_1;
wire na2445_1_i;
wire na2446_2;
wire na2446_2_i;
wire na2447_1;
wire na2447_1_i;
wire na2448_2;
wire na2448_2_i;
wire na2449_1;
wire na2449_1_i;
wire na2450_2;
wire na2450_2_i;
wire na2451_1;
wire na2451_1_i;
wire na2451_2;
wire na2451_2_i;
wire na2452_1;
wire na2452_1_i;
wire na2453_2;
wire na2453_2_i;
wire na2454_1;
wire na2454_1_i;
wire na2455_2;
wire na2455_2_i;
wire na2456_1;
wire na2456_1_i;
wire na2456_2;
wire na2456_2_i;
wire na2457_1;
wire na2457_1_i;
wire na2458_2;
wire na2458_2_i;
wire na2459_1;
wire na2459_1_i;
wire na2460_2;
wire na2460_2_i;
wire na2461_1;
wire na2461_1_i;
wire na2462_2;
wire na2462_2_i;
wire na2463_1;
wire na2463_1_i;
wire na2464_1;
wire na2464_1_i;
wire na2464_2;
wire na2464_2_i;
wire na2465_2;
wire na2465_2_i;
wire na2466_1;
wire na2466_1_i;
wire na2467_1;
wire na2467_1_i;
wire na2467_2;
wire na2467_2_i;
wire na2468_2;
wire na2468_2_i;
wire na2469_1;
wire na2469_1_i;
wire na2470_2;
wire na2470_2_i;
wire na2471_1;
wire na2471_1_i;
wire na2471_2;
wire na2471_2_i;
wire na2472_1;
wire na2472_1_i;
wire na2473_1;
wire na2473_1_i;
wire na2474_1;
wire na2474_1_i;
wire na2474_2;
wire na2474_2_i;
wire na2475_1;
wire na2475_1_i;
wire na2475_2;
wire na2475_2_i;
wire na2476_1;
wire na2476_1_i;
wire na2477_2;
wire na2477_2_i;
wire na2478_1;
wire na2478_1_i;
wire na2479_2;
wire na2479_2_i;
wire na2480_1;
wire na2480_1_i;
wire na2480_2;
wire na2480_2_i;
wire na2481_1;
wire na2481_1_i;
wire na2482_2;
wire na2482_2_i;
wire na2483_1;
wire na2483_1_i;
wire na2484_2;
wire na2484_2_i;
wire na2485_1;
wire na2485_1_i;
wire na2486_2;
wire na2486_2_i;
wire na2487_1;
wire na2487_1_i;
wire na2488_2;
wire na2488_2_i;
wire na2489_1;
wire na2489_1_i;
wire na2490_2;
wire na2490_2_i;
wire na2491_1;
wire na2491_1_i;
wire na2492_2;
wire na2492_2_i;
wire na2493_1;
wire na2493_1_i;
wire na2494_2;
wire na2494_2_i;
wire na2495_1;
wire na2495_1_i;
wire na2496_2;
wire na2496_2_i;
wire na2497_1;
wire na2497_1_i;
wire na2498_2;
wire na2498_2_i;
wire na2499_1;
wire na2499_1_i;
wire na2500_2;
wire na2500_2_i;
wire na2501_1;
wire na2501_1_i;
wire na2502_2;
wire na2502_2_i;
wire na2503_1;
wire na2503_1_i;
wire na2504_2;
wire na2504_2_i;
wire na2505_2;
wire na2505_2_i;
wire na2506_2;
wire na2506_2_i;
wire na2507_1;
wire na2507_1_i;
wire na2508_2;
wire na2508_2_i;
wire na2509_1;
wire na2509_1_i;
wire na2510_2;
wire na2510_2_i;
wire na2511_1;
wire na2511_1_i;
wire na2512_2;
wire na2512_2_i;
wire na2513_1;
wire na2513_1_i;
wire na2514_2;
wire na2514_2_i;
wire na2515_1;
wire na2515_1_i;
wire na2516_2;
wire na2516_2_i;
wire na2517_1;
wire na2517_1_i;
wire na2518_2;
wire na2518_2_i;
wire na2519_1;
wire na2519_1_i;
wire na2520_2;
wire na2520_2_i;
wire na2521_1;
wire na2521_1_i;
wire na2522_2;
wire na2522_2_i;
wire na2523_1;
wire na2523_1_i;
wire na2524_2;
wire na2524_2_i;
wire na2525_1;
wire na2525_1_i;
wire na2526_2;
wire na2526_2_i;
wire na2527_1;
wire na2527_1_i;
wire na2528_2;
wire na2528_2_i;
wire na2529_1;
wire na2529_1_i;
wire na2530_2;
wire na2530_2_i;
wire na2531_1;
wire na2531_1_i;
wire na2532_2;
wire na2532_2_i;
wire na2533_1;
wire na2533_1_i;
wire na2534_2;
wire na2534_2_i;
wire na2535_2;
wire na2535_2_i;
wire na2536_2;
wire na2536_2_i;
wire na2537_1;
wire na2537_1_i;
wire na2538_2;
wire na2538_2_i;
wire na2539_1;
wire na2539_1_i;
wire na2540_2;
wire na2540_2_i;
wire na2541_1;
wire na2541_1_i;
wire na2542_2;
wire na2542_2_i;
wire na2543_1;
wire na2543_1_i;
wire na2544_2;
wire na2544_2_i;
wire na2545_1;
wire na2545_1_i;
wire na2546_2;
wire na2546_2_i;
wire na2547_1;
wire na2547_1_i;
wire na2548_2;
wire na2548_2_i;
wire na2549_1;
wire na2549_1_i;
wire na2550_2;
wire na2550_2_i;
wire na2551_1;
wire na2551_1_i;
wire na2552_2;
wire na2552_2_i;
wire na2553_1;
wire na2553_1_i;
wire na2554_2;
wire na2554_2_i;
wire na2555_1;
wire na2555_1_i;
wire na2556_2;
wire na2556_2_i;
wire na2557_1;
wire na2557_1_i;
wire na2558_2;
wire na2558_2_i;
wire na2559_1;
wire na2559_1_i;
wire na2560_2;
wire na2560_2_i;
wire na2561_1;
wire na2561_1_i;
wire na2562_2;
wire na2562_2_i;
wire na2563_1;
wire na2563_1_i;
wire na2564_1;
wire na2564_1_i;
wire na2565_1;
wire na2565_1_i;
wire na2566_2;
wire na2566_2_i;
wire na2567_1;
wire na2567_1_i;
wire na2568_2;
wire na2568_2_i;
wire na2569_1;
wire na2569_1_i;
wire na2570_2;
wire na2570_2_i;
wire na2571_1;
wire na2571_1_i;
wire na2572_2;
wire na2572_2_i;
wire na2573_1;
wire na2573_1_i;
wire na2574_2;
wire na2574_2_i;
wire na2575_1;
wire na2575_1_i;
wire na2576_2;
wire na2576_2_i;
wire na2577_1;
wire na2577_1_i;
wire na2578_2;
wire na2578_2_i;
wire na2579_1;
wire na2579_1_i;
wire na2580_2;
wire na2580_2_i;
wire na2581_1;
wire na2581_1_i;
wire na2582_2;
wire na2582_2_i;
wire na2583_1;
wire na2583_1_i;
wire na2584_2;
wire na2584_2_i;
wire na2585_1;
wire na2585_1_i;
wire na2586_2;
wire na2586_2_i;
wire na2587_1;
wire na2587_1_i;
wire na2588_2;
wire na2588_2_i;
wire na2589_1;
wire na2589_1_i;
wire na2590_2;
wire na2590_2_i;
wire na2591_1;
wire na2591_1_i;
wire na2592_2;
wire na2592_2_i;
wire na2593_1;
wire na2593_1_i;
wire na2594_1;
wire na2594_1_i;
wire na2595_1;
wire na2595_1_i;
wire na2596_2;
wire na2596_2_i;
wire na2597_1;
wire na2597_1_i;
wire na2598_2;
wire na2598_2_i;
wire na2599_1;
wire na2599_1_i;
wire na2600_2;
wire na2600_2_i;
wire na2601_1;
wire na2601_1_i;
wire na2602_2;
wire na2602_2_i;
wire na2603_1;
wire na2603_1_i;
wire na2604_2;
wire na2604_2_i;
wire na2605_1;
wire na2605_1_i;
wire na2606_2;
wire na2606_2_i;
wire na2607_1;
wire na2607_1_i;
wire na2608_2;
wire na2608_2_i;
wire na2609_1;
wire na2609_1_i;
wire na2610_2;
wire na2610_2_i;
wire na2611_1;
wire na2611_1_i;
wire na2612_2;
wire na2612_2_i;
wire na2613_1;
wire na2613_1_i;
wire na2614_2;
wire na2614_2_i;
wire na2615_1;
wire na2615_1_i;
wire na2616_2;
wire na2616_2_i;
wire na2617_1;
wire na2617_1_i;
wire na2618_2;
wire na2618_2_i;
wire na2619_1;
wire na2619_1_i;
wire na2620_2;
wire na2620_2_i;
wire na2621_1;
wire na2621_1_i;
wire na2622_2;
wire na2622_2_i;
wire na2623_2;
wire na2623_2_i;
wire na2624_2;
wire na2624_2_i;
wire na2625_1;
wire na2625_1_i;
wire na2626_2;
wire na2626_2_i;
wire na2627_1;
wire na2627_1_i;
wire na2628_2;
wire na2628_2_i;
wire na2629_1;
wire na2629_1_i;
wire na2630_2;
wire na2630_2_i;
wire na2631_1;
wire na2631_1_i;
wire na2632_2;
wire na2632_2_i;
wire na2633_1;
wire na2633_1_i;
wire na2634_2;
wire na2634_2_i;
wire na2635_1;
wire na2635_1_i;
wire na2636_2;
wire na2636_2_i;
wire na2637_1;
wire na2637_1_i;
wire na2638_2;
wire na2638_2_i;
wire na2639_1;
wire na2639_1_i;
wire na2640_2;
wire na2640_2_i;
wire na2641_1;
wire na2641_1_i;
wire na2642_2;
wire na2642_2_i;
wire na2643_1;
wire na2643_1_i;
wire na2644_2;
wire na2644_2_i;
wire na2645_1;
wire na2645_1_i;
wire na2646_2;
wire na2646_2_i;
wire na2647_1;
wire na2647_1_i;
wire na2648_2;
wire na2648_2_i;
wire na2649_1;
wire na2649_1_i;
wire na2650_2;
wire na2650_2_i;
wire na2651_1;
wire na2651_1_i;
wire na2652_2;
wire na2652_2_i;
wire na2653_2;
wire na2653_2_i;
wire na2654_2;
wire na2654_2_i;
wire na2655_1;
wire na2655_1_i;
wire na2656_2;
wire na2656_2_i;
wire na2657_1;
wire na2657_1_i;
wire na2658_2;
wire na2658_2_i;
wire na2659_1;
wire na2659_1_i;
wire na2660_2;
wire na2660_2_i;
wire na2661_1;
wire na2661_1_i;
wire na2662_2;
wire na2662_2_i;
wire na2663_1;
wire na2663_1_i;
wire na2664_2;
wire na2664_2_i;
wire na2665_1;
wire na2665_1_i;
wire na2666_2;
wire na2666_2_i;
wire na2667_1;
wire na2667_1_i;
wire na2668_2;
wire na2668_2_i;
wire na2669_1;
wire na2669_1_i;
wire na2670_2;
wire na2670_2_i;
wire na2671_1;
wire na2671_1_i;
wire na2672_2;
wire na2672_2_i;
wire na2673_1;
wire na2673_1_i;
wire na2674_2;
wire na2674_2_i;
wire na2675_1;
wire na2675_1_i;
wire na2676_2;
wire na2676_2_i;
wire na2677_1;
wire na2677_1_i;
wire na2678_2;
wire na2678_2_i;
wire na2679_1;
wire na2679_1_i;
wire na2680_2;
wire na2680_2_i;
wire na2681_1;
wire na2681_1_i;
wire na2682_1;
wire na2682_1_i;
wire na2683_1;
wire na2683_1_i;
wire na2684_2;
wire na2684_2_i;
wire na2685_1;
wire na2685_1_i;
wire na2686_2;
wire na2686_2_i;
wire na2687_1;
wire na2687_1_i;
wire na2688_2;
wire na2688_2_i;
wire na2689_1;
wire na2689_1_i;
wire na2690_2;
wire na2690_2_i;
wire na2691_1;
wire na2691_1_i;
wire na2692_2;
wire na2692_2_i;
wire na2693_1;
wire na2693_1_i;
wire na2694_2;
wire na2694_2_i;
wire na2695_1;
wire na2695_1_i;
wire na2696_2;
wire na2696_2_i;
wire na2697_1;
wire na2697_1_i;
wire na2698_2;
wire na2698_2_i;
wire na2699_1;
wire na2699_1_i;
wire na2700_2;
wire na2700_2_i;
wire na2701_1;
wire na2701_1_i;
wire na2702_2;
wire na2702_2_i;
wire na2703_1;
wire na2703_1_i;
wire na2704_2;
wire na2704_2_i;
wire na2705_1;
wire na2705_1_i;
wire na2706_2;
wire na2706_2_i;
wire na2707_1;
wire na2707_1_i;
wire na2708_2;
wire na2708_2_i;
wire na2709_1;
wire na2709_1_i;
wire na2710_2;
wire na2710_2_i;
wire na2711_2;
wire na2711_2_i;
wire na2712_2;
wire na2712_2_i;
wire na2713_1;
wire na2713_1_i;
wire na2714_2;
wire na2714_2_i;
wire na2715_1;
wire na2715_1_i;
wire na2716_2;
wire na2716_2_i;
wire na2717_1;
wire na2717_1_i;
wire na2718_2;
wire na2718_2_i;
wire na2719_1;
wire na2719_1_i;
wire na2720_2;
wire na2720_2_i;
wire na2721_1;
wire na2721_1_i;
wire na2722_2;
wire na2722_2_i;
wire na2723_1;
wire na2723_1_i;
wire na2724_2;
wire na2724_2_i;
wire na2725_1;
wire na2725_1_i;
wire na2726_2;
wire na2726_2_i;
wire na2727_1;
wire na2727_1_i;
wire na2728_2;
wire na2728_2_i;
wire na2729_1;
wire na2729_1_i;
wire na2730_2;
wire na2730_2_i;
wire na2731_1;
wire na2731_1_i;
wire na2732_2;
wire na2732_2_i;
wire na2733_1;
wire na2733_1_i;
wire na2734_2;
wire na2734_2_i;
wire na2735_1;
wire na2735_1_i;
wire na2736_2;
wire na2736_2_i;
wire na2737_1;
wire na2737_1_i;
wire na2738_2;
wire na2738_2_i;
wire na2739_1;
wire na2739_1_i;
wire na2740_1;
wire na2740_1_i;
wire na2741_1;
wire na2741_1_i;
wire na2742_2;
wire na2742_2_i;
wire na2743_1;
wire na2743_1_i;
wire na2745_2;
wire na2745_2_i;
wire na2746_1;
wire na2746_1_i;
wire na2748_2;
wire na2748_2_i;
wire na2749_1;
wire na2749_1_i;
wire na2750_2;
wire na2750_2_i;
wire na2752_1;
wire na2752_1_i;
wire na2753_2;
wire na2753_2_i;
wire na2756_1;
wire na2756_1_i;
wire na2757_2;
wire na2757_2_i;
wire na2758_1;
wire na2758_1_i;
wire na2759_2;
wire na2759_2_i;
wire na2761_1;
wire na2761_1_i;
wire na2762_2;
wire na2762_2_i;
wire na2763_1;
wire na2763_1_i;
wire na2764_2;
wire na2764_2_i;
wire na2765_1;
wire na2765_1_i;
wire na2766_2;
wire na2766_2_i;
wire na2767_1;
wire na2767_1_i;
wire na2768_2;
wire na2768_2_i;
wire na2769_1;
wire na2769_1_i;
wire na2770_2;
wire na2770_2_i;
wire na2771_1;
wire na2771_1_i;
wire na2772_2;
wire na2772_2_i;
wire na2773_1;
wire na2773_1_i;
wire na2774_2;
wire na2774_2_i;
wire na2775_1;
wire na2775_1_i;
wire na2776_1;
wire na2776_1_i;
wire na2777_1;
wire na2777_1_i;
wire na2778_2;
wire na2778_2_i;
wire na2779_1;
wire na2779_1_i;
wire na2780_2;
wire na2780_2_i;
wire na2781_1;
wire na2781_1_i;
wire na2782_2;
wire na2782_2_i;
wire na2783_1;
wire na2783_1_i;
wire na2784_2;
wire na2784_2_i;
wire na2785_1;
wire na2785_1_i;
wire na2786_2;
wire na2786_2_i;
wire na2787_1;
wire na2787_1_i;
wire na2788_2;
wire na2788_2_i;
wire na2789_1;
wire na2789_1_i;
wire na2790_2;
wire na2790_2_i;
wire na2791_1;
wire na2791_1_i;
wire na2792_2;
wire na2792_2_i;
wire na2793_1;
wire na2793_1_i;
wire na2794_2;
wire na2794_2_i;
wire na2795_1;
wire na2795_1_i;
wire na2796_2;
wire na2796_2_i;
wire na2797_1;
wire na2797_1_i;
wire na2798_2;
wire na2798_2_i;
wire na2799_1;
wire na2799_1_i;
wire na2800_2;
wire na2800_2_i;
wire na2801_1;
wire na2801_1_i;
wire na2802_2;
wire na2802_2_i;
wire na2803_1;
wire na2803_1_i;
wire na2804_2;
wire na2804_2_i;
wire na2805_2;
wire na2805_2_i;
wire na2806_2;
wire na2806_2_i;
wire na2807_1;
wire na2807_1_i;
wire na2808_2;
wire na2808_2_i;
wire na2809_1;
wire na2809_1_i;
wire na2810_2;
wire na2810_2_i;
wire na2811_1;
wire na2811_1_i;
wire na2812_2;
wire na2812_2_i;
wire na2813_1;
wire na2813_1_i;
wire na2814_2;
wire na2814_2_i;
wire na2815_1;
wire na2815_1_i;
wire na2816_2;
wire na2816_2_i;
wire na2817_1;
wire na2817_1_i;
wire na2818_2;
wire na2818_2_i;
wire na2819_1;
wire na2819_1_i;
wire na2820_2;
wire na2820_2_i;
wire na2821_1;
wire na2821_1_i;
wire na2822_2;
wire na2822_2_i;
wire na2823_1;
wire na2823_1_i;
wire na2824_2;
wire na2824_2_i;
wire na2825_1;
wire na2825_1_i;
wire na2826_2;
wire na2826_2_i;
wire na2827_1;
wire na2827_1_i;
wire na2828_2;
wire na2828_2_i;
wire na2829_1;
wire na2829_1_i;
wire na2830_2;
wire na2830_2_i;
wire na2831_1;
wire na2831_1_i;
wire na2832_2;
wire na2832_2_i;
wire na2833_1;
wire na2833_1_i;
wire na2834_2;
wire na2834_2_i;
wire na2835_2;
wire na2835_2_i;
wire na2836_2;
wire na2836_2_i;
wire na2837_1;
wire na2837_1_i;
wire na2838_2;
wire na2838_2_i;
wire na2839_1;
wire na2839_1_i;
wire na2841_2;
wire na2841_2_i;
wire na2842_1;
wire na2842_1_i;
wire na2844_2;
wire na2844_2_i;
wire na2845_1;
wire na2845_1_i;
wire na2846_2;
wire na2846_2_i;
wire na2848_1;
wire na2848_1_i;
wire na2849_2;
wire na2849_2_i;
wire na2852_1;
wire na2852_1_i;
wire na2853_2;
wire na2853_2_i;
wire na2854_1;
wire na2854_1_i;
wire na2855_2;
wire na2855_2_i;
wire na2857_1;
wire na2857_1_i;
wire na2858_2;
wire na2858_2_i;
wire na2860_1;
wire na2860_1_i;
wire na2861_2;
wire na2861_2_i;
wire na2862_1;
wire na2862_1_i;
wire na2863_2;
wire na2863_2_i;
wire na2865_1;
wire na2865_1_i;
wire na2866_2;
wire na2866_2_i;
wire na2867_1;
wire na2867_1_i;
wire na2868_2;
wire na2868_2_i;
wire na2869_1;
wire na2869_1_i;
wire na2870_2;
wire na2870_2_i;
wire na2871_1;
wire na2871_1_i;
wire na2872_1;
wire na2872_1_i;
wire na2873_1;
wire na2873_1_i;
wire na2874_2;
wire na2874_2_i;
wire na2875_1;
wire na2875_1_i;
wire na2876_2;
wire na2876_2_i;
wire na2877_1;
wire na2877_1_i;
wire na2878_2;
wire na2878_2_i;
wire na2879_1;
wire na2879_1_i;
wire na2880_2;
wire na2880_2_i;
wire na2881_1;
wire na2881_1_i;
wire na2882_2;
wire na2882_2_i;
wire na2883_1;
wire na2883_1_i;
wire na2884_2;
wire na2884_2_i;
wire na2885_1;
wire na2885_1_i;
wire na2886_2;
wire na2886_2_i;
wire na2887_1;
wire na2887_1_i;
wire na2888_2;
wire na2888_2_i;
wire na2889_1;
wire na2889_1_i;
wire na2890_2;
wire na2890_2_i;
wire na2891_1;
wire na2891_1_i;
wire na2892_2;
wire na2892_2_i;
wire na2893_1;
wire na2893_1_i;
wire na2894_2;
wire na2894_2_i;
wire na2895_1;
wire na2895_1_i;
wire na2896_2;
wire na2896_2_i;
wire na2897_1;
wire na2897_1_i;
wire na2898_2;
wire na2898_2_i;
wire na2899_1;
wire na2899_1_i;
wire na2900_2;
wire na2900_2_i;
wire na2901_1;
wire na2901_1_i;
wire na2902_1;
wire na2902_1_i;
wire na2903_1;
wire na2903_1_i;
wire na2904_2;
wire na2904_2_i;
wire na2905_1;
wire na2905_1_i;
wire na2906_2;
wire na2906_2_i;
wire na2907_1;
wire na2907_1_i;
wire na2908_2;
wire na2908_2_i;
wire na2909_1;
wire na2909_1_i;
wire na2910_2;
wire na2910_2_i;
wire na2911_1;
wire na2911_1_i;
wire na2912_2;
wire na2912_2_i;
wire na2913_1;
wire na2913_1_i;
wire na2914_2;
wire na2914_2_i;
wire na2915_1;
wire na2915_1_i;
wire na2916_2;
wire na2916_2_i;
wire na2917_1;
wire na2917_1_i;
wire na2918_2;
wire na2918_2_i;
wire na2919_1;
wire na2919_1_i;
wire na2920_2;
wire na2920_2_i;
wire na2921_1;
wire na2921_1_i;
wire na2922_2;
wire na2922_2_i;
wire na2923_1;
wire na2923_1_i;
wire na2924_2;
wire na2924_2_i;
wire na2925_1;
wire na2925_1_i;
wire na2926_2;
wire na2926_2_i;
wire na2927_1;
wire na2927_1_i;
wire na2928_2;
wire na2928_2_i;
wire na2929_1;
wire na2929_1_i;
wire na2930_2;
wire na2930_2_i;
wire na2931_2;
wire na2931_2_i;
wire na2932_2;
wire na2932_2_i;
wire na2933_1;
wire na2933_1_i;
wire na2934_2;
wire na2934_2_i;
wire na2935_1;
wire na2935_1_i;
wire na2936_2;
wire na2936_2_i;
wire na2937_1;
wire na2937_1_i;
wire na2938_2;
wire na2938_2_i;
wire na2939_1;
wire na2939_1_i;
wire na2940_2;
wire na2940_2_i;
wire na2941_1;
wire na2941_1_i;
wire na2942_2;
wire na2942_2_i;
wire na2943_1;
wire na2943_1_i;
wire na2944_2;
wire na2944_2_i;
wire na2945_1;
wire na2945_1_i;
wire na2946_1;
wire na2946_1_i;
wire na2946_2;
wire na2946_2_i;
wire na2949_1;
wire na2949_1_i;
wire na2949_2;
wire na2949_2_i;
wire na2950_2;
wire na2950_2_i;
wire na2953_1;
wire na2953_1_i;
wire na2953_2;
wire na2953_2_i;
wire na2955_1;
wire na2955_1_i;
wire na2956_1;
wire na2956_1_i;
wire na2956_2;
wire na2956_2_i;
wire na2957_1;
wire na2957_1_i;
wire na2957_2;
wire na2957_2_i;
wire na2959_1;
wire na2959_1_i;
wire na2959_2;
wire na2959_2_i;
wire na2961_1;
wire na2961_1_i;
wire na2961_2;
wire na2961_2_i;
wire na2963_2;
wire na2963_2_i;
wire na2964_1;
wire na2964_1_i;
wire na2965_1;
wire na2965_1_i;
wire na2965_2;
wire na2965_2_i;
wire na2966_1;
wire na2966_1_i;
wire na2966_2;
wire na2966_2_i;
wire na2967_1;
wire na2967_1_i;
wire na2967_2;
wire na2967_2_i;
wire na2968_1;
wire na2968_1_i;
wire na2968_2;
wire na2968_2_i;
wire na2969_1;
wire na2969_1_i;
wire na2969_2;
wire na2969_2_i;
wire na2970_2;
wire na2970_2_i;
wire na2971_1;
wire na2971_1_i;
wire na2976_1;
wire na2976_1_i;
wire na2976_2;
wire na2976_2_i;
wire na2978_2;
wire na2978_2_i;
wire na2979_1;
wire na2979_1_i;
wire na2980_2;
wire na2980_2_i;
wire na2981_1;
wire na2981_1_i;
wire na2982_2;
wire na2982_2_i;
wire na2983_1;
wire na2983_1_i;
wire na2984_2;
wire na2984_2_i;
wire na2985_1;
wire na2985_1_i;
wire na2986_2;
wire na2986_2_i;
wire na2987_2;
wire na2987_2_i;
wire na2988_2;
wire na2988_2_i;
wire na2989_1;
wire na2989_1_i;
wire na2990_2;
wire na2990_2_i;
wire na2991_1;
wire na2991_1_i;
wire na2992_2;
wire na2992_2_i;
wire na2993_1;
wire na2993_1_i;
wire na2994_2;
wire na2994_2_i;
wire na2995_1;
wire na2995_1_i;
wire na2996_2;
wire na2996_2_i;
wire na2997_1;
wire na2997_1_i;
wire na2998_2;
wire na2998_2_i;
wire na2999_1;
wire na2999_1_i;
wire na3000_2;
wire na3000_2_i;
wire na3001_1;
wire na3001_1_i;
wire na3002_2;
wire na3002_2_i;
wire na3003_1;
wire na3003_1_i;
wire na3004_2;
wire na3004_2_i;
wire na3005_1;
wire na3005_1_i;
wire na3006_2;
wire na3006_2_i;
wire na3007_1;
wire na3007_1_i;
wire na3008_2;
wire na3008_2_i;
wire na3009_1;
wire na3009_1_i;
wire na3010_2;
wire na3010_2_i;
wire na3011_1;
wire na3011_1_i;
wire na3013_2;
wire na3013_2_i;
wire na3014_1;
wire na3014_1_i;
wire na3015_2;
wire na3015_2_i;
wire na3016_1;
wire na3016_1_i;
wire na3017_1;
wire na3017_1_i;
wire na3017_2;
wire na3017_2_i;
wire na3018_1;
wire na3018_1_i;
wire na3019_1;
wire na3019_1_i;
wire na3021_2;
wire na3021_2_i;
wire na3022_1;
wire na3022_1_i;
wire na3023_2;
wire na3023_2_i;
wire na3024_1;
wire na3024_1_i;
wire na3025_1;
wire na3025_1_i;
wire na3025_2;
wire na3025_2_i;
wire na3026_2;
wire na3026_2_i;
wire na3027_1;
wire na3027_1_i;
wire na3029_2;
wire na3029_2_i;
wire na3030_1;
wire na3030_1_i;
wire na3031_2;
wire na3031_2_i;
wire na3032_1;
wire na3032_1_i;
wire na3033_1;
wire na3033_1_i;
wire na3033_2;
wire na3033_2_i;
wire na3034_2;
wire na3034_2_i;
wire na3035_1;
wire na3035_1_i;
wire na3037_2;
wire na3037_2_i;
wire na3038_1;
wire na3038_1_i;
wire na3039_2;
wire na3039_2_i;
wire na3040_1;
wire na3040_1_i;
wire na3041_1;
wire na3041_1_i;
wire na3041_2;
wire na3041_2_i;
wire na3042_2;
wire na3042_2_i;
wire na3043_1;
wire na3043_1_i;
wire na3044_2;
wire na3044_2_i;
wire na3045_1;
wire na3045_1_i;
wire na3046_2;
wire na3046_2_i;
wire na3047_1;
wire na3047_1_i;
wire na3048_2;
wire na3048_2_i;
wire na3049_1;
wire na3049_1_i;
wire na3050_2;
wire na3050_2_i;
wire na3051_1;
wire na3051_1_i;
wire na3052_2;
wire na3052_2_i;
wire na3053_1;
wire na3053_1_i;
wire na3054_1;
wire na3054_1_i;
wire na3055_1;
wire na3055_1_i;
wire na3056_2;
wire na3056_2_i;
wire na3057_1;
wire na3057_1_i;
wire na3058_2;
wire na3058_2_i;
wire na3059_1;
wire na3059_1_i;
wire na3060_2;
wire na3060_2_i;
wire na3061_1;
wire na3061_1_i;
wire na3062_2;
wire na3062_2_i;
wire na3063_1;
wire na3063_1_i;
wire na3064_2;
wire na3064_2_i;
wire na3065_1;
wire na3065_1_i;
wire na3066_2;
wire na3066_2_i;
wire na3067_1;
wire na3067_1_i;
wire na3068_2;
wire na3068_2_i;
wire na3069_1;
wire na3069_1_i;
wire na3070_2;
wire na3070_2_i;
wire na3071_1;
wire na3071_1_i;
wire na3072_2;
wire na3072_2_i;
wire na3073_1;
wire na3073_1_i;
wire na3074_2;
wire na3074_2_i;
wire na3075_1;
wire na3075_1_i;
wire na3076_2;
wire na3076_2_i;
wire na3077_1;
wire na3077_1_i;
wire na3078_2;
wire na3078_2_i;
wire na3079_1;
wire na3079_1_i;
wire na3080_2;
wire na3080_2_i;
wire na3081_1;
wire na3081_1_i;
wire na3082_2;
wire na3082_2_i;
wire na3083_2;
wire na3083_2_i;
wire na3084_2;
wire na3084_2_i;
wire na3085_1;
wire na3085_1_i;
wire na3086_2;
wire na3086_2_i;
wire na3087_1;
wire na3087_1_i;
wire na3088_2;
wire na3088_2_i;
wire na3089_1;
wire na3089_1_i;
wire na3090_2;
wire na3090_2_i;
wire na3091_1;
wire na3091_1_i;
wire na3092_2;
wire na3092_2_i;
wire na3093_1;
wire na3093_1_i;
wire na3094_2;
wire na3094_2_i;
wire na3095_1;
wire na3095_1_i;
wire na3096_2;
wire na3096_2_i;
wire na3097_1;
wire na3097_1_i;
wire na3098_2;
wire na3098_2_i;
wire na3099_1;
wire na3099_1_i;
wire na3100_2;
wire na3100_2_i;
wire na3101_1;
wire na3101_1_i;
wire na3102_2;
wire na3102_2_i;
wire na3103_1;
wire na3103_1_i;
wire na3104_2;
wire na3104_2_i;
wire na3105_1;
wire na3105_1_i;
wire na3106_2;
wire na3106_2_i;
wire na3107_1;
wire na3107_1_i;
wire na3108_2;
wire na3108_2_i;
wire na3109_1;
wire na3109_1_i;
wire na3110_2;
wire na3110_2_i;
wire na3111_1;
wire na3111_1_i;
wire na3112_2;
wire na3112_2_i;
wire na3113_2;
wire na3113_2_i;
wire na3114_2;
wire na3114_2_i;
wire na3115_1;
wire na3115_1_i;
wire na3116_2;
wire na3116_2_i;
wire na3117_1;
wire na3117_1_i;
wire na3118_2;
wire na3118_2_i;
wire na3119_1;
wire na3119_1_i;
wire na3120_2;
wire na3120_2_i;
wire na3121_1;
wire na3121_1_i;
wire na3122_2;
wire na3122_2_i;
wire na3123_1;
wire na3123_1_i;
wire na3124_2;
wire na3124_2_i;
wire na3125_1;
wire na3125_1_i;
wire na3126_2;
wire na3126_2_i;
wire na3127_1;
wire na3127_1_i;
wire na3128_2;
wire na3128_2_i;
wire na3129_1;
wire na3129_1_i;
wire na3130_2;
wire na3130_2_i;
wire na3131_1;
wire na3131_1_i;
wire na3132_2;
wire na3132_2_i;
wire na3133_1;
wire na3133_1_i;
wire na3134_2;
wire na3134_2_i;
wire na3135_1;
wire na3135_1_i;
wire na3136_2;
wire na3136_2_i;
wire na3137_1;
wire na3137_1_i;
wire na3138_2;
wire na3138_2_i;
wire na3139_1;
wire na3139_1_i;
wire na3140_2;
wire na3140_2_i;
wire na3141_1;
wire na3141_1_i;
wire na3142_1;
wire na3142_1_i;
wire na3143_1;
wire na3143_1_i;
wire na3144_2;
wire na3144_2_i;
wire na3145_1;
wire na3145_1_i;
wire na3146_2;
wire na3146_2_i;
wire na3147_1;
wire na3147_1_i;
wire na3148_2;
wire na3148_2_i;
wire na3149_1;
wire na3149_1_i;
wire na3150_2;
wire na3150_2_i;
wire na3151_1;
wire na3151_1_i;
wire na3151_2;
wire na3151_2_i;
wire na3153_1;
wire na3153_1_i;
wire na3154_2;
wire na3154_2_i;
wire na3155_1;
wire na3155_1_i;
wire na3156_2;
wire na3156_2_i;
wire na3157_1;
wire na3157_1_i;
wire na3158_2;
wire na3158_2_i;
wire na3159_1;
wire na3159_1_i;
wire na3160_2;
wire na3160_2_i;
wire na3161_1;
wire na3161_1_i;
wire na3162_2;
wire na3162_2_i;
wire na3163_1;
wire na3163_1_i;
wire na3164_2;
wire na3164_2_i;
wire na3165_1;
wire na3165_1_i;
wire na3166_2;
wire na3166_2_i;
wire na3167_1;
wire na3167_1_i;
wire na3168_2;
wire na3168_2_i;
wire na3169_1;
wire na3169_1_i;
wire na3170_1;
wire na3170_1_i;
wire na3170_2;
wire na3170_2_i;
wire na3172_2;
wire na3172_2_i;
wire na3173_1;
wire na3173_1_i;
wire na3174_2;
wire na3174_2_i;
wire na3175_1;
wire na3175_1_i;
wire na3175_2;
wire na3175_2_i;
wire na3176_1;
wire na3176_1_i;
wire na3178_1;
wire na3178_1_i;
wire na3180_1;
wire na3180_1_i;
wire na3181_1;
wire na3181_1_i;
wire na3181_2;
wire na3181_2_i;
wire na3182_1;
wire na3182_1_i;
wire na3182_2;
wire na3182_2_i;
wire na3184_2;
wire na3184_2_i;
wire na3185_1;
wire na3185_1_i;
wire na3186_2;
wire na3186_2_i;
wire na3187_1;
wire na3187_1_i;
wire na3188_2;
wire na3188_2_i;
wire na3189_1;
wire na3189_1_i;
wire na3190_2;
wire na3190_2_i;
wire na3191_1;
wire na3191_1_i;
wire na3192_2;
wire na3192_2_i;
wire na3193_1;
wire na3193_1_i;
wire na3194_2;
wire na3194_2_i;
wire na3195_1;
wire na3195_1_i;
wire na3196_2;
wire na3196_2_i;
wire na3197_1;
wire na3197_1_i;
wire na3198_2;
wire na3198_2_i;
wire na3199_1;
wire na3199_1_i;
wire na3200_2;
wire na3200_2_i;
wire na3201_1;
wire na3201_1_i;
wire na3202_2;
wire na3202_2_i;
wire na3203_1;
wire na3203_1_i;
wire na3204_2;
wire na3204_2_i;
wire na3205_1;
wire na3205_1_i;
wire na3206_2;
wire na3206_2_i;
wire na3207_1;
wire na3207_1_i;
wire na3208_2;
wire na3208_2_i;
wire na3209_1;
wire na3209_1_i;
wire na3210_2;
wire na3210_2_i;
wire na3211_2;
wire na3211_2_i;
wire na3212_2;
wire na3212_2_i;
wire na3213_1;
wire na3213_1_i;
wire na3214_1;
wire na3214_1_i;
wire na3214_2;
wire na3214_2_i;
wire na3215_2;
wire na3215_2_i;
wire na3216_1;
wire na3216_1_i;
wire na3216_2;
wire na3216_2_i;
wire na3217_1;
wire na3217_1_i;
wire na3219_2;
wire na3219_2_i;
wire na3220_1;
wire na3220_1_i;
wire na3220_2;
wire na3220_2_i;
wire na3223_1;
wire na3223_1_i;
wire na3223_2;
wire na3223_2_i;
wire na3225_1;
wire na3225_1_i;
wire na3226_2;
wire na3226_2_i;
wire na3227_1;
wire na3227_1_i;
wire na3228_2;
wire na3228_2_i;
wire na3229_1;
wire na3229_1_i;
wire na3230_2;
wire na3230_2_i;
wire na3231_1;
wire na3231_1_i;
wire na3232_2;
wire na3232_2_i;
wire na3234_1;
wire na3234_1_i;
wire na3235_1;
wire na3235_1_i;
wire na3235_2;
wire na3235_2_i;
wire na3236_1;
wire na3237_1;
wire na3238_1;
wire na3239_1;
wire na3240_1;
wire na3241_1;
wire na3242_1;
wire na3243_1;
wire na3244_1;
wire na3245_1;
wire na3246_1;
wire na3247_1;
wire na3248_1;
wire na3249_1;
wire na3250_1;
wire na3251_1;
wire na3252_1;
wire na3253_1;
wire na3254_1;
wire na3255_1;
wire na3256_1;
wire na3257_1;
wire na3258_1;
wire na3259_1;
wire na3260_1;
wire na3261_1;
wire na3262_1;
wire na3263_1;
wire na3264_1;
wire na3265_1;
wire na3266_1;
wire na3267_1;
wire na3268_1;
wire na3269_1;
wire na3277_1;
wire na3278_1;
wire na3278_2;
wire na3280_1;
wire na3280_4;
wire na3281_1;
wire na3283_2;
wire na3284_1;
wire na3285_2;
wire na3286_1;
wire na3286_2;
wire na3289_1;
wire na3290_2;
wire na3291_1;
wire na3291_2;
wire na3294_1;
wire na3295_1;
wire na3296_1;
wire na3296_2;
wire na3299_2;
wire na3300_2;
wire na3301_1;
wire na3301_2;
wire na3304_2;
wire na3305_1;
wire na3306_1;
wire na3306_2;
wire na3309_2;
wire na3310_2;
wire na3311_1;
wire na3311_2;
wire na3314_1;
wire na3315_2;
wire na3316_1;
wire na3316_2;
wire na3319_1;
wire na3320_1;
wire na3321_1;
wire na3321_2;
wire na3324_2;
wire na3325_1;
wire na3326_1;
wire na3326_2;
wire na3329_2;
wire na3330_1;
wire na3331_1;
wire na3331_2;
wire na3334_2;
wire na3335_2;
wire na3336_1;
wire na3336_2;
wire na3339_2;
wire na3340_1;
wire na3341_1;
wire na3341_2;
wire na3344_2;
wire na3345_2;
wire na3347_1;
wire na3349_2;
wire na3350_1;
wire na3351_1;
wire na3351_2;
wire na3354_1;
wire na3355_2;
wire na3356_1;
wire na3356_2;
wire na3359_1;
wire na3360_2;
wire na3361_1;
wire na3361_2;
wire na3364_1;
wire na3365_1;
wire na3366_1;
wire na3366_2;
wire na3369_1;
wire na3370_1;
wire na3371_1;
wire na3371_2;
wire na3374_2;
wire na3375_1;
wire na3376_1;
wire na3376_2;
wire na3379_2;
wire na3380_1;
wire na3381_1;
wire na3381_2;
wire na3384_2;
wire na3385_1;
wire na3386_1;
wire na3386_2;
wire na3389_2;
wire na3390_2;
wire na3391_1;
wire na3391_2;
wire na3394_1;
wire na3395_1;
wire na3397_1;
wire na3399_2;
wire na3400_1;
wire na3401_1;
wire na3401_2;
wire na3404_1;
wire na3405_2;
wire na3406_1;
wire na3406_2;
wire na3409_2;
wire na3410_1;
wire na3411_1;
wire na3411_2;
wire na3414_2;
wire na3415_2;
wire na3416_1;
wire na3416_2;
wire na3419_2;
wire na3420_1;
wire na3421_1;
wire na3421_2;
wire na3424_2;
wire na3425_2;
wire na3426_1;
wire na3426_2;
wire na3429_2;
wire na3430_1;
wire na3431_1;
wire na3431_2;
wire na3434_2;
wire na3435_1;
wire na3436_1;
wire na3436_2;
wire na3439_1;
wire na3440_2;
wire na3441_1;
wire na3442_2;
wire na3446_1;
wire na3447_1;
wire na3449_2;
wire na3451_1;
wire na3452_2;
wire na3453_1;
wire na3454_2;
wire na3455_1;
wire na3456_2;
wire na3457_2;
wire na3462_1;
wire na3463_2;
wire na3465_1;
wire na3466_1;
wire na3470_1;
wire na3472_2;
wire na3474_1;
wire na3475_2;
wire na3479_1;
wire na3480_2;
wire na3483_2;
wire na3484_1;
wire na3486_1;
wire na3489_1;
wire na3490_2;
wire na3492_2;
wire na3494_1;
wire na3495_2;
wire na3499_1;
wire na3502_1;
wire na3503_1;
wire na3505_2;
wire na3507_2;
wire na3508_1;
wire na3512_1;
wire na3513_2;
wire na3516_1;
wire na3518_2;
wire na3519_1;
wire na3519_2;
wire na3523_1;
wire na3528_1;
wire na3528_2;
wire na3529_1;
wire na3531_1;
wire na3532_1;
wire na3533_2;
wire na3534_1;
wire na3534_2;
wire na3540_1;
wire na3541_1;
wire na3542_1;
wire na3543_1;
wire na3543_2;
wire na3548_2;
wire na3550_2;
wire na3551_1;
wire na3551_2;
wire na3555_1;
wire na3556_1;
wire na3557_2;
wire na3558_1;
wire na3558_2;
wire na3563_1;
wire na3565_1;
wire na3566_1;
wire na3566_2;
wire na3570_1;
wire na3570_2;
wire na3572_1;
wire na3576_1;
wire na3577_2;
wire na3579_1;
wire na3580_1;
wire na3580_2;
wire na3585_1;
wire na3585_2;
wire na3590_2;
wire na3592_1;
wire na3593_1;
wire na3593_2;
wire na3597_2;
wire na3598_1;
wire na3599_1;
wire na3599_2;
wire na3604_2;
wire na3606_1;
wire na3607_1;
wire na3607_2;
wire na3611_1;
wire na3612_1;
wire na3614_2;
wire na3615_1;
wire na3615_2;
wire na3620_1;
wire na3621_2;
wire na3622_1;
wire na3622_2;
wire na3627_1;
wire na3627_2;
wire na3629_1;
wire na3633_1;
wire na3634_1;
wire na3635_2;
wire na3636_1;
wire na3636_2;
wire na3641_1;
wire na3642_1;
wire na3643_2;
wire na3644_1;
wire na3644_2;
wire na3650_1;
wire na3651_1;
wire na3652_2;
wire na3653_1;
wire na3653_2;
wire na3659_1;
wire na3663_1;
wire na3663_2;
wire na3665_1;
wire na3667_2;
wire na3668_1;
wire na3668_2;
wire na3672_1;
wire na3673_1;
wire na3674_1;
wire na3675_1;
wire na3675_2;
wire na3680_1;
wire na3681_2;
wire na3682_1;
wire na3683_1;
wire na3683_2;
wire na3689_1;
wire na3689_2;
wire na3694_2;
wire na3695_1;
wire na3696_1;
wire na3699_2;
wire na3700_1;
wire na3704_2;
wire na3705_1;
wire na3707_2;
wire na3709_1;
wire na3711_1;
wire na3712_2;
wire na3713_1;
wire na3714_2;
wire na3716_1;
wire na3717_1;
wire na3717_2;
wire na3720_1;
wire na3721_1;
wire na3722_2;
wire na3723_1;
wire na3724_1;
wire na3726_2;
wire na3728_2;
wire na3729_2;
wire na3730_1;
wire na3731_2;
wire na3732_1;
wire na3733_1;
wire na3734_2;
wire na3735_1;
wire na3736_2;
wire na3737_1;
wire na3738_2;
wire na3739_1;
wire na3741_2;
wire na3742_1;
wire na3744_2;
wire na3748_2;
wire na3749_1;
wire na3750_2;
wire na3751_1;
wire na3752_2;
wire na3756_1;
wire na3757_2;
wire na3758_1;
wire na3759_2;
wire na3760_1;
wire na3761_2;
wire na3762_2;
wire na3764_1;
wire na3766_2;
wire na3767_2;
wire na3768_1;
wire na3769_2;
wire na3770_2;
wire na3771_1;
wire na3772_1;
wire na3773_2;
wire na3774_2;
wire na3775_1;
wire na3778_2;
wire na3781_1;
wire na3782_2;
wire na3784_1;
wire na3785_2;
wire na3788_2;
wire na3790_1;
wire na3792_2;
wire na3794_1;
wire na3795_1;
wire na3796_2;
wire na3798_1;
wire na3799_2;
wire na3800_1;
wire na3801_2;
wire na3803_1;
wire na3805_2;
wire na3806_1;
wire na3807_2;
wire na3808_1;
wire na3809_2;
wire na3810_1;
wire na3811_2;
wire na3812_1;
wire na3813_2;
wire na3814_1;
wire na3863_2;
wire na3864_1;
wire na3865_2;
wire na3866_1;
wire na3867_2;
wire na3868_1;
wire na3869_1;
wire na3870_2;
wire na3944_1;
wire na3945_1;
wire na3946_2;
wire na3947_1;
wire na3948_1;
wire na3950_1;
wire na3951_1;
wire na3952_1;
wire na3953_2;
wire na3954_2;
wire na3955_1;
wire na3956_2;
wire na3957_1;
wire na3958_1;
wire na3959_1;
wire na3959_2;
wire na3960_2;
wire na3962_1;
wire na3963_1;
wire na3964_2;
wire na3965_1;
wire na3966_2;
wire na3975_1;
wire na3975_2;
wire na3976_2;
wire na3978_2;
wire na3979_1;
wire na3980_1;
wire na3981_2;
wire na3983_1;
wire na3984_1;
wire na3984_2;
wire na3990_1;
wire na3990_2;
wire na3991_1;
wire na3993_1;
wire na3994_1;
wire na3995_2;
wire na3996_1;
wire na3997_2;
wire na4006_1;
wire na4006_2;
wire na4007_2;
wire na4009_1;
wire na4010_1;
wire na4011_1;
wire na4012_1;
wire na4013_1;
wire na4014_1;
wire na4015_2;
wire na4018_1;
wire na4019_2;
wire na4020_1;
wire na4021_2;
wire na4022_1;
wire na4023_2;
wire na4024_1;
wire na4025_2;
wire na4026_1;
wire na4027_2;
wire na4028_1;
wire na4029_2;
wire na4030_1;
wire na4031_2;
wire na4034_1;
wire na4035_2;
wire na4036_2;
wire na4037_1;
wire na4038_2;
wire na4039_1;
wire na4040_2;
wire na4041_1;
wire na4042_1;
wire na4043_2;
wire na4044_1;
wire na4045_1;
wire na4054_1;
wire na4054_2;
wire na4055_1;
wire na4057_2;
wire na4058_1;
wire na4059_1;
wire na4059_2;
wire na4060_1;
wire na4061_1;
wire na4061_2;
wire na4063_2;
wire na4066_1;
wire na4067_2;
wire na4068_1;
wire na4068_2;
wire na4071_1;
wire na4072_2;
wire na4073_2;
wire na4076_2;
wire na4079_1;
wire na4082_1;
wire na4083_1;
wire na4085_1;
wire na4088_2;
wire na4089_1;
wire na4093_1;
wire na4100_2;
wire na4101_1;
wire na4102_2;
wire na4103_1;
wire na4104_1;
wire na4105_2;
wire na4107_1;
wire na4109_2;
wire na4110_1;
wire na4111_2;
wire na4112_1;
wire na4114_1;
wire na4115_1;
wire na4116_1;
wire na4117_1;
wire na4119_1;
wire na4120_1;
wire na4121_2;
wire na4122_1;
wire na4124_2;
wire na4125_1;
wire na4126_2;
wire na4127_1;
wire na4129_2;
wire na4130_1;
wire na4131_2;
wire na4132_1;
wire na4134_2;
wire na4135_1;
wire na4136_1;
wire na4141_2;
wire na4146_1;
wire na4147_1;
wire na4151_1;
wire na4152_2;
wire na4153_1;
wire na4154_2;
wire na4155_2;
wire na4156_2;
wire na4157_2;
wire na4158_2;
wire na4159_2;
wire na4160_2;
wire na4161_2;
wire na4162_2;
wire na4163_2;
wire na4164_2;
wire na4165_2;
wire na4166_2;
wire na4167_2;
wire na4168_2;
wire na4169_2;
wire na4170_2;
wire na4171_2;
wire na4172_2;
wire na4173_2;
wire na4174_2;
wire na4175_2;
wire na4176_2;
wire na4177_2;
wire na4178_2;
wire na4179_2;
wire na4180_2;
wire na4181_2;
wire na4182_2;
wire na4183_2;
wire na4184_2;
wire na4185_2;
wire na4186_2;
wire na4187_2;
wire na4188_2;
wire na4189_2;
wire na4190_2;
wire na4191_2;
wire na4192_2;
wire na4193_2;
wire na4194_2;
wire na4195_2;
wire na4196_2;
wire na4197_2;
wire na4198_2;
wire na4199_2;
wire na4200_2;
wire na4201_2;
wire na4202_2;
wire na4203_2;
wire na4204_2;
wire na4205_2;
wire na4206_2;
wire na4207_2;
wire na4208_2;
wire na4209_2;
wire na4210_2;
wire na4211_2;
wire na4212_2;
wire na4213_2;
wire na4214_2;
wire na4215_2;
wire na4216_2;
wire na4217_2;
wire na4218_2;
wire na4219_2;
wire na4220_2;
wire na4221_2;
wire na4222_2;
wire na4223_2;
wire na4224_2;
wire na4225_2;
wire na4226_2;
wire na4227_2;
wire na4228_2;
wire na4229_2;
wire na4230_2;
wire na4231_2;
wire na4232_2;
wire na4233_2;
wire na4234_2;
wire na4235_2;
wire na4236_2;
wire na4237_2;
wire na4238_2;
wire na4239_2;
wire na4240_2;
wire na4241_2;
wire na4242_2;
wire na4243_2;
wire na4244_2;
wire na4245_2;
wire na4246_2;
wire na4247_2;
wire na4248_2;
wire na4249_2;
wire na4250_2;
wire na4251_2;
wire na4252_2;
wire na4253_2;
wire na4254_2;
wire na4255_2;
wire na4256_2;
wire na4257_2;
wire na4258_2;
wire na4259_2;
wire na4260_2;
wire na4261_2;
wire na4262_2;
wire na4263_2;
wire na4264_2;
wire na4265_2;
wire na4266_2;
wire na4267_2;
wire na4268_2;
wire na4269_2;
wire na4270_2;
wire na4271_2;
wire na4272_2;
wire na4273_2;
wire na4274_2;
wire na4275_2;
wire na4276_2;
wire na4277_2;
wire na4278_2;
wire na4279_2;
wire na4280_2;
wire na4281_2;
wire na4282_2;
wire na4283_2;
wire na4284_2;
wire na4285_2;
wire na4286_2;
wire na4287_2;
wire na4288_2;
wire na4289_2;
wire na4290_2;
wire na4291_2;
wire na4292_2;
wire na4293_2;
wire na4294_2;
wire na4295_2;
wire na4296_2;
wire na4297_2;
wire na4298_2;
wire na4299_2;
wire na4300_2;
wire na4301_2;
wire na4302_2;
wire na4303_2;
wire na4304_2;
wire na4305_2;
wire na4306_2;
wire na4307_2;
wire na4308_2;
wire na4309_2;
wire na4310_2;
wire na4311_2;
wire na4312_2;
wire na4313_2;
wire na4314_2;
wire na4315_2;
wire na4316_2;
wire na4317_2;
wire na4318_2;
wire na4319_2;
wire na4320_2;
wire na4321_2;
wire na4322_2;
wire na4323_2;
wire na4324_2;
wire na4325_2;
wire na4326_2;
wire na4327_2;
wire na4328_2;
wire na4329_2;
wire na4330_2;
wire na4331_2;
wire na4332_2;
wire na4333_2;
wire na4334_2;
wire na4335_2;
wire na4336_2;
wire na4337_2;
wire na4338_2;
wire na4339_2;
wire na4340_2;
wire na4341_2;
wire na4342_2;
wire na4343_2;
wire na4344_2;
wire na4345_2;
wire na4346_2;
wire na4347_2;
wire na4348_2;
wire na4349_2;
wire na4350_2;
wire na4351_2;
wire na4352_2;
wire na4353_2;
wire na4354_2;
wire na4355_2;
wire na4356_2;
wire na4357_2;
wire na4358_2;
wire na4359_2;
wire na4360_2;
wire na4361_2;
wire na4362_2;
wire na4363_2;
wire na4364_2;
wire na4365_2;
wire na4366_2;
wire na4367_2;
wire na4368_2;
wire na4369_2;
wire na4370_2;
wire na4371_2;
wire na4372_2;
wire na4373_2;
wire na4374_2;
wire na4375_2;
wire na4376_2;
wire na4377_2;
wire na4378_2;
wire na4379_2;
wire na4380_2;
wire na4381_2;
wire na4382_2;
wire na4383_2;
wire na4384_2;
wire na4385_2;
wire na4386_2;
wire na4387_2;
wire na4388_2;
wire na4389_2;
wire na4390_2;
wire na4391_2;
wire na4392_2;
wire na4393_2;
wire na4394_2;
wire na4395_2;
wire na4396_2;
wire na4397_2;
wire na4398_2;
wire na4399_2;
wire na4400_2;
wire na4401_2;
wire na4402_2;
wire na4403_2;
wire na4404_2;
wire na4405_2;
wire na4406_2;
wire na4407_2;
wire na4408_2;
wire na4409_2;
wire na4410_2;
wire na4411_2;
wire na4412_2;
wire na4413_2;
wire na4414_2;
wire na4415_2;
wire na4416_2;
wire na4481_1;
wire na4481_2;
wire na4481_3;
wire na4481_6;
wire na4154_10;
wire na4155_10;
wire na4156_10;
wire na4157_10;
wire na4158_10;
wire na4159_10;
wire na4160_10;

// C_AND////      x87y104     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_2), .IN6(1'b1), .IN7(na3169_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y108     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1860_1), .IN7(na3169_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y110     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3_4 ( .OUT(na3_2), .IN1(1'b1), .IN2(na1860_2), .IN3(na3169_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y112     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1862_1), .IN6(1'b1), .IN7(na3169_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y112     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2), .IN1(na1862_2), .IN2(1'b1), .IN3(na3169_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y115     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1864_1), .IN7(na3169_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y85     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7_4 ( .OUT(na7_2), .IN1(1'b1), .IN2(~na1957_2), .IN3(na1958_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y86     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4161_2), .IN7(~na1930_2), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y83     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2), .IN1(na1866_1), .IN2(1'b1), .IN3(na7_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y87     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1866_2), .IN6(1'b1), .IN7(na7_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x149y85     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a11_4 ( .OUT(na11_2), .IN1(1'b1), .IN2(na1868_1), .IN3(na7_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y88     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1868_2), .IN7(na7_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x98y97     80'h00_0018_00_0000_0EEE_E0EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(na22_2), .IN2(1'b0), .IN3(na20_1), .IN4(na18_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3278_1), .IN8(na4395_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a14 ( .PCLK0(na14_1), .PCLK1(_d0), .PCLK2(_d1), .PCLK3(_d2), .CLK0(na3268_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0), .SER_CLK(1'b0),
                  .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_///AND/      x127y81     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a15_4 ( .OUT(na15_2), .IN1(1'b1), .IN2(na16_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y82     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a16_4 ( .OUT(na16_2), .IN1(1'b1), .IN2(1'b1), .IN3(na17_1), .IN4(~na3150_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y71     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4382_2), .IN6(1'b1), .IN7(na3151_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y102     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na4336_2), .IN8(na2279_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x110y96     80'h00_0018_00_0000_0CEE_BA00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4382_2), .IN6(1'b0), .IN7(na3151_1), .IN8(~na3150_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x106y97     80'h00_0018_00_0040_0C05_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1), .IN1(na2458_2), .IN2(1'b0), .IN3(na2418_2), .IN4(1'b0), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na4310_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x123y83     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a21_4 ( .OUT(na21_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na17_1), .IN4(~na3150_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x97y95     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a22_4 ( .OUT(na22_2), .IN1(~na25_1), .IN2(na3283_2), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y93     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2416_2), .IN7(1'b1), .IN8(~na24_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y90     80'h00_0060_00_0000_0C08_FF51
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a24_4 ( .OUT(na24_2), .IN1(~na2415_2), .IN2(~na2416_1), .IN3(~na2417_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y95     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2834_2), .IN8(~na3284_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y83     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a26_4 ( .OUT(na26_2), .IN1(1'b1), .IN2(~na3285_2), .IN3(~na3151_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y84     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na16_2), .IN7(1'b1), .IN8(na4310_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x110y98     80'h00_0018_00_0000_0EEE_ACCE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1), .IN1(na31_1), .IN2(na3286_2), .IN3(1'b0), .IN4(na30_1), .IN5(1'b0), .IN6(na3286_1), .IN7(na32_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y98     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(na2459_1), .IN6(na4312_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y99     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2771_1), .IN6(na2280_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x110y95     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a32_4 ( .OUT(na32_2), .IN1(na3289_1), .IN2(~na33_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y98     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2835_2), .IN8(~na3290_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x108y79     80'h00_0018_00_0000_0EEE_CCEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_1 ( .OUT(na34_1), .IN1(1'b0), .IN2(na3291_2), .IN3(na38_1), .IN4(na36_1), .IN5(1'b0), .IN6(na3291_1), .IN7(1'b0), .IN8(na39_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y82     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na37_1), .IN6(na3294_1), .IN7(~na26_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y79     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2836_2), .IN6(1'b0), .IN7(~na3295_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y75     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2772_2), .IN8(na2281_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y84     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2420_2), .IN6(1'b0), .IN7(na2460_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x100y96     80'h00_0018_00_0000_0EEE_0EEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a40_1 ( .OUT(na40_1), .IN1(1'b0), .IN2(na3296_2), .IN3(na42_1), .IN4(na43_1), .IN5(na44_2), .IN6(na3296_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y105     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2282_2), .IN6(na2773_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y102     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(~na4165_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2461_1),
                    .IN8(na4314_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x99y101     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a44_4 ( .OUT(na44_2), .IN1(~na45_1), .IN2(na3299_2), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y99     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2837_1), .IN6(~na3300_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y71     80'h00_0018_00_0000_0EEE_CCAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1), .IN1(na50_1), .IN2(na3301_2), .IN3(na48_1), .IN4(1'b0), .IN5(1'b0), .IN6(na3301_1), .IN7(1'b0), .IN8(na51_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y83     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3304_2), .IN6(~na49_1), .IN7(~na26_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y88     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3305_1), .IN8(~na2838_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y87     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2283_2), .IN6(na4337_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y84     80'h00_0018_00_0040_0A50_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(na2462_2), .IN6(1'b0), .IN7(na4315_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x104y77     80'h00_0018_00_0000_0EEE_ACEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a52_1 ( .OUT(na52_1), .IN1(na55_1), .IN2(1'b0), .IN3(na3306_2), .IN4(na54_1), .IN5(1'b0), .IN6(na56_2), .IN7(na3306_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y82     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(na2463_1), .IN6(na2423_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y83     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2775_1), .IN6(na2284_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x105y72     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a56_4 ( .OUT(na56_2), .IN1(na3309_2), .IN2(~na58_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x105y70     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a57_4 ( .OUT(na57_2), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y82     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3310_2), .IN8(~na2839_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x104y86     80'h00_0018_00_0000_0EEE_CCEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1), .IN1(na62_1), .IN2(1'b0), .IN3(na61_1), .IN4(na3311_2), .IN5(1'b0), .IN6(na63_2), .IN7(1'b0), .IN8(na3311_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y87     80'h00_0018_00_0040_0AA0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(na2464_1), .IN7(1'b0), .IN8(na2424_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y89     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2776_1), .IN8(na2285_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x103y84     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a63_4 ( .OUT(na63_2), .IN1(na3314_1), .IN2(~na64_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y90     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3315_2), .IN6(~na2464_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y69     80'h00_0018_00_0000_0EEE_CCEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1), .IN1(na69_1), .IN2(1'b0), .IN3(na67_1), .IN4(na3316_2), .IN5(1'b0), .IN6(na70_1), .IN7(1'b0), .IN8(na3316_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x108y71     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3319_1), .IN6(~na68_1), .IN7(~na26_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y72     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_1 ( .OUT(na68_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3320_1), .IN6(~na2841_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y77     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2286_2), .IN8(na2777_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y76     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2425_2), .IN6(1'b0), .IN7(na2465_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x122y98     80'h00_0018_00_0000_0EEE_ACCE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a71_1 ( .OUT(na71_1), .IN1(na73_2), .IN2(na3321_2), .IN3(1'b0), .IN4(na75_1), .IN5(1'b0), .IN6(na3321_1), .IN7(na76_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x119y103     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a73_4 ( .OUT(na73_2), .IN1(na3324_2), .IN2(~na74_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y102     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na3325_1), .IN7(1'b0), .IN8(~na2842_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y108     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2778_2), .IN6(na4306_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y103     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na4165_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2426_1), .IN8(na2466_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x134y98     80'h00_0018_00_0000_0EEE_E0CE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a77_1 ( .OUT(na77_1), .IN1(na81_1), .IN2(na79_2), .IN3(1'b0), .IN4(na3326_2), .IN5(1'b0), .IN6(1'b0), .IN7(na82_1), .IN8(na3326_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x127y94     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a79_4 ( .OUT(na79_2), .IN1(na3329_2), .IN2(~na80_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y98     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3330_1), .IN6(~na2467_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y99     80'h00_0018_00_0040_0AA0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(1'b1), .IN2(~na4164_2), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(na2779_1), .IN7(1'b0), .IN8(na2288_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y95     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a82_1 ( .OUT(na82_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na4165_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2427_1), .IN8(na4329_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x127y97     80'h00_0018_00_0000_0EEE_CE0E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1), .IN1(na86_1), .IN2(na3331_2), .IN3(1'b0), .IN4(1'b0), .IN5(na85_1), .IN6(na3331_1), .IN7(1'b0), .IN8(na87_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y95     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(~na4165_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4330_2),
                    .IN8(na2428_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y99     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2780_2), .IN6(na2289_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x120y96     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3334_2), .IN6(~na88_1), .IN7(~na26_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y98     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3335_2), .IN6(~na2844_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x111y105     80'h00_0018_00_0000_0EEE_0EEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1), .IN1(na3336_2), .IN2(1'b0), .IN3(na92_1), .IN4(na91_1), .IN5(na3336_1), .IN6(na93_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y106     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a91_1 ( .OUT(na91_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2781_1), .IN6(na2290_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y103     80'h00_0018_00_0040_0AA0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(na2469_1), .IN7(1'b0), .IN8(na2429_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x113y102     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3339_2), .IN6(~na94_1), .IN7(~na26_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y100     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2845_1), .IN6(1'b0), .IN7(~na3340_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x122y87     80'h00_0018_00_0000_0EEE_0EEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a95_1 ( .OUT(na95_1), .IN1(na3341_2), .IN2(1'b0), .IN3(na97_1), .IN4(na98_1), .IN5(na3341_1), .IN6(na99_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y91     80'h00_0018_00_0040_0A50_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(na4331_2), .IN6(1'b0), .IN7(na2430_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y94     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_1 ( .OUT(na98_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2291_1), .IN6(na2782_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x119y90     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na100_1), .IN6(na3344_2), .IN7(~na26_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y93     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2846_2), .IN6(~na3345_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x109y76     80'h00_0018_00_0000_0888_3BE5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a101_1 ( .OUT(na101_1), .IN1(~na106_1), .IN2(1'b0), .IN3(na26_2), .IN4(na3347_1), .IN5(na3350_1), .IN6(~na16_2), .IN7(1'b0),
                     .IN8(~na105_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y78     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3349_2), .IN6(~na2471_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y78     80'h00_0018_00_0040_0AA0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(na2471_1), .IN7(1'b0), .IN8(na2431_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y79     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2783_1), .IN8(na4307_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x115y94     80'h00_0018_00_0000_0EEE_CAAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1), .IN1(na3351_2), .IN2(na110_1), .IN3(na109_1), .IN4(1'b0), .IN5(na3351_1), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na111_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y97     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a109_1 ( .OUT(na109_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na4338_2), .IN8(na2293_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y94     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2432_1), .IN6(1'b0), .IN7(na2472_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x112y92     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a111_4 ( .OUT(na111_2), .IN1(na3354_1), .IN2(~na112_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y96     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2848_1), .IN6(1'b0), .IN7(~na3355_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x94y79     80'h00_0018_00_0000_0EEE_CCEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1), .IN1(na117_1), .IN2(1'b0), .IN3(na115_2), .IN4(na3356_2), .IN5(1'b0), .IN6(na118_1), .IN7(1'b0),
                     .IN8(na3356_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x104y69     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a115_4 ( .OUT(na115_2), .IN1(na3359_1), .IN2(~na116_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x99y78     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a116_1 ( .OUT(na116_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3360_2), .IN8(~na2849_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y77     80'h00_0018_00_0040_0A50_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b1), .IN2(na4164_2), .IN3(1'b1), .IN4(na4310_2), .IN5(na2785_1), .IN6(1'b0), .IN7(na2294_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y76     80'h00_0018_00_0040_0A50_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(na2473_1), .IN6(1'b0), .IN7(na2433_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x132y102     80'h00_0018_00_0000_0EEE_CCAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1), .IN1(na123_1), .IN2(na3361_2), .IN3(na121_2), .IN4(1'b0), .IN5(1'b0), .IN6(na3361_1), .IN7(1'b0),
                     .IN8(na124_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x122y95     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a121_4 ( .OUT(na121_2), .IN1(na3364_1), .IN2(~na122_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y98     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2474_2), .IN6(1'b0), .IN7(~na3365_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y97     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(na2474_1), .IN6(na2434_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y100     80'h00_0018_00_0040_0A50_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a124_1 ( .OUT(na124_1), .IN1(1'b1), .IN2(na4164_2), .IN3(1'b1), .IN4(na4310_2), .IN5(na2786_2), .IN6(1'b0), .IN7(na2295_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x139y95     80'h00_0018_00_0000_0EEE_ECCC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1), .IN1(1'b0), .IN2(na129_1), .IN3(1'b0), .IN4(na3366_2), .IN5(1'b0), .IN6(na127_1), .IN7(na130_1),
                     .IN8(na3366_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x125y94     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na128_1), .IN6(na3369_1), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y95     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2475_2), .IN8(~na3370_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y98     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a129_1 ( .OUT(na129_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na4308_2), .IN6(na2787_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y93     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a130_1 ( .OUT(na130_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2435_1), .IN6(1'b0), .IN7(na2475_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x120y102     80'h00_0018_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_1 ( .OUT(na131_1), .IN1(1'b0), .IN2(na133_1), .IN3(na3371_2), .IN4(na135_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3371_1),
                     .IN8(na136_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x115y96     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3374_2), .IN6(~na134_1), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y98     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2852_1), .IN6(1'b0), .IN7(~na3375_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y104     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a135_1 ( .OUT(na135_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2788_2), .IN6(na2297_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y98     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(~na4165_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2476_1),
                     .IN8(na2436_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x122y96     80'h00_0018_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a137_1 ( .OUT(na137_1), .IN1(na139_1), .IN2(na141_1), .IN3(na3376_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3376_1),
                     .IN8(na142_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x115y97     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a139_1 ( .OUT(na139_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3379_2), .IN6(~na140_1), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x115y100     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(~na2853_2), .IN2(~na3380_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2416_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y106     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2789_1), .IN8(na2298_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y100     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2437_1), .IN6(1'b0), .IN7(na2477_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x117y86     80'h00_0018_00_0000_0EEE_ACCE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a143_1 ( .OUT(na143_1), .IN1(na145_2), .IN2(na3381_2), .IN3(1'b0), .IN4(na147_1), .IN5(1'b0), .IN6(na3381_1), .IN7(na148_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x115y85     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a145_4 ( .OUT(na145_2), .IN1(~na146_1), .IN2(na3384_2), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y87     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3385_1), .IN6(~na2854_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y90     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a147_1 ( .OUT(na147_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(na2478_1), .IN6(na4318_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y91     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2299_1), .IN6(na2790_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x110y66     80'h00_0018_00_0000_0EEE_ECAC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a149_1 ( .OUT(na149_1), .IN1(1'b0), .IN2(na151_2), .IN3(na3386_2), .IN4(1'b0), .IN5(1'b0), .IN6(na153_1), .IN7(na3386_1),
                     .IN8(na154_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x105y68     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a151_4 ( .OUT(na151_2), .IN1(~na152_1), .IN2(na3389_2), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y75     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(~na2855_2), .IN7(1'b0), .IN8(~na3390_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y76     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a153_1 ( .OUT(na153_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2300_2), .IN6(na2791_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y74     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1), .IN1(1'b1), .IN2(na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(na2439_2), .IN6(na2479_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x120y79     80'h00_0018_00_0000_0EEE_CAEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b0), .IN2(na157_1), .IN3(na158_1), .IN4(na3391_2), .IN5(na159_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na3391_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y84     80'h00_0018_00_0040_0A50_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(na2480_1), .IN6(1'b0), .IN7(na2440_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y85     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a158_1 ( .OUT(na158_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2792_2), .IN6(na2301_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x117y85     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a159_4 ( .OUT(na159_2), .IN1(~na160_1), .IN2(na3394_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y87     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_1 ( .OUT(na160_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2480_2), .IN6(~na3395_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x109y84     80'h00_0018_00_0000_0888_5BE5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(~na166_1), .IN2(1'b0), .IN3(na26_2), .IN4(na3397_1), .IN5(na3400_1), .IN6(~na16_2), .IN7(~na165_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y81     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a163_1 ( .OUT(na163_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na3399_2), .IN7(1'b0), .IN8(~na2857_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y85     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_1 ( .OUT(na165_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na4339_2), .IN6(na2302_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y83     80'h00_0018_00_0040_0A50_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(na2481_1), .IN6(1'b0), .IN7(na2441_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x106y98     80'h00_0018_00_0000_0EEE_CCEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_1 ( .OUT(na167_1), .IN1(na169_1), .IN2(1'b0), .IN3(na170_1), .IN4(na3401_2), .IN5(1'b0), .IN6(na171_1), .IN7(1'b0),
                     .IN8(na3401_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y97     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a169_1 ( .OUT(na169_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(na2450_2), .IN6(na2442_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y105     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_1 ( .OUT(na170_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2303_1), .IN8(na2794_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x103y100     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a171_1 ( .OUT(na171_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na172_1), .IN6(na3404_1), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y103     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a172_1 ( .OUT(na172_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(~na2858_2), .IN7(1'b0), .IN8(~na3405_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x129y99     80'h00_0018_00_0000_0EEE_AAEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(1'b0), .IN2(na177_1), .IN3(na3406_2), .IN4(na175_1), .IN5(na178_1), .IN6(1'b0), .IN7(na3406_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x120y98     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a175_1 ( .OUT(na175_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3409_2), .IN6(~na176_1), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y100     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a176_1 ( .OUT(na176_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4310_2), .IN5(~na3410_1), .IN6(1'b0), .IN7(~na2451_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y98     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2443_1), .IN6(1'b0), .IN7(na2451_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y97     80'h00_0018_00_0040_0AA0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(1'b1), .IN2(~na4164_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(na2304_2), .IN7(1'b0),
                     .IN8(na2795_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x118y107     80'h00_0018_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b0), .IN2(na182_1), .IN3(na3411_2), .IN4(na181_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3411_1),
                     .IN8(na183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y104     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2305_1), .IN6(na2796_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y104     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2444_2), .IN6(1'b0), .IN7(na2452_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x116y104     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na184_1), .IN6(na3414_2), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y103     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a184_1 ( .OUT(na184_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2860_1), .IN6(1'b0), .IN7(~na3415_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x106y100     80'h00_0018_00_0000_0EEE_AAEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a185_1 ( .OUT(na185_1), .IN1(1'b0), .IN2(na188_1), .IN3(na3416_2), .IN4(na187_1), .IN5(na189_2), .IN6(1'b0), .IN7(na3416_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y102     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a187_1 ( .OUT(na187_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(na2445_1), .IN6(1'b0), .IN7(na4323_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y106     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na4340_2), .IN6(na2306_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x115y97     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a189_4 ( .OUT(na189_2), .IN1(na3419_2), .IN2(~na190_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y100     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a190_1 ( .OUT(na190_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na3420_1), .IN7(1'b0), .IN8(~na2861_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y96     80'h00_0018_00_0000_0EEE_0ECE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a191_1 ( .OUT(na191_1), .IN1(na3421_2), .IN2(na193_2), .IN3(1'b0), .IN4(na195_1), .IN5(na3421_1), .IN6(na196_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x105y92     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a193_4 ( .OUT(na193_2), .IN1(na3424_2), .IN2(~na194_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y98     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2862_1), .IN6(1'b0), .IN7(~na3425_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y100     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a195_1 ( .OUT(na195_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2798_2), .IN6(na2307_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y96     80'h00_0018_00_0040_0AA0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a196_1 ( .OUT(na196_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(na2446_2), .IN7(1'b0), .IN8(na2454_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x104y88     80'h00_0018_00_0000_0EEE_ECAA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a197_1 ( .OUT(na197_1), .IN1(na199_1), .IN2(1'b0), .IN3(na3426_2), .IN4(1'b0), .IN5(1'b0), .IN6(na200_1), .IN7(na3426_1),
                     .IN8(na201_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y87     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(~na4165_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2455_2),
                     .IN8(na2447_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y94     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a200_1 ( .OUT(na200_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2799_1), .IN6(na2308_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x104y82     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a201_4 ( .OUT(na201_2), .IN1(na3429_2), .IN2(~na202_1), .IN3(~na26_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y88     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2863_2), .IN6(1'b0), .IN7(~na3430_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x109y92     80'h00_0018_00_0000_0EEE_0EEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a203_1 ( .OUT(na203_1), .IN1(1'b0), .IN2(na3431_2), .IN3(na207_1), .IN4(na205_1), .IN5(na208_1), .IN6(na3431_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x104y94     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a205_1 ( .OUT(na205_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na206_1), .IN6(na3434_2), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y91     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a206_1 ( .OUT(na206_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(~na2456_2), .IN7(1'b0), .IN8(~na3435_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y97     80'h00_0018_00_0040_0A50_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(1'b1), .IN2(na4164_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(na2309_1), .IN6(1'b0), .IN7(na2800_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y93     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_1 ( .OUT(na208_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na4165_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2448_2),
                     .IN8(na4324_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x108y89     80'h00_0018_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a209_1 ( .OUT(na209_1), .IN1(1'b0), .IN2(na211_1), .IN3(na213_1), .IN4(na3436_2), .IN5(1'b0), .IN6(1'b0), .IN7(na214_1),
                     .IN8(na3436_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x105y92     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a211_1 ( .OUT(na211_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3439_1), .IN6(~na212_1), .IN7(~na26_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y92     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2865_1), .IN6(1'b0), .IN7(~na3440_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y93     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a213_1 ( .OUT(na213_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2310_2), .IN6(na4341_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y87     80'h00_0018_00_0040_0AA0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(na2457_1), .IN7(1'b0), .IN8(na4321_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x118y99     80'h00_0060_00_0000_0C06_FF65
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a215_4 ( .OUT(na215_2), .IN1(~na4174_2), .IN2(1'b0), .IN3(na259_1), .IN4(na258_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x120y104     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a216_4 ( .OUT(na216_2), .IN1(~na255_2), .IN2(na249_1), .IN3(na4175_2), .IN4(~na256_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y103     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a217_1 ( .OUT(na217_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na218_1), .IN6(1'b0), .IN7(na243_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y109     80'h00_0018_00_0040_0A72_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1), .IN1(na219_1), .IN2(1'b1), .IN3(1'b1), .IN4(na239_1), .IN5(na3441_1), .IN6(~na241_1), .IN7(na240_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y111     80'h00_0018_00_0040_0AF1_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a219_1 ( .OUT(na219_1), .IN1(1'b1), .IN2(~na232_1), .IN3(~na1799_1), .IN4(1'b1), .IN5(~na3442_2), .IN6(na1797_1), .IN7(na4396_2),
                     .IN8(na1801_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y113     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a220_4 ( .OUT(na220_2), .IN1(na3017_2), .IN2(na3013_2), .IN3(~na3015_2), .IN4(~na4358_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y114     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a221_4 ( .OUT(na221_2), .IN1(na3017_1), .IN2(1'b0), .IN3(~na3011_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x124y113     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a222_4 ( .OUT(na222_2), .IN1(~na3016_1), .IN2(na3014_1), .IN3(na3011_1), .IN4(na4358_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x125y113     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a223_1 ( .OUT(na223_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3016_1), .IN6(na3014_1), .IN7(na3015_2), .IN8(~na4356_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y118     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na236_1), .IN8(~na230_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y116     80'h00_0018_00_0040_0AD2_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_1 ( .OUT(na225_1), .IN1(na226_1), .IN2(1'b1), .IN3(~na222_2), .IN4(1'b1), .IN5(na3010_2), .IN6(1'b1), .IN7(na3446_1),
                     .IN8(na227_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y113     80'h00_0018_00_0000_0C66_A900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3016_1), .IN6(na3014_1), .IN7(na3015_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x128y114     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3017_2), .IN6(na3014_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x125y115     80'h00_0060_00_0000_0C08_FF56
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a228_4 ( .OUT(na228_2), .IN1(~na223_1), .IN2(na4180_2), .IN3(na222_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y110     80'h00_0018_00_0040_0A98_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(na3017_2), .IN2(1'b1), .IN3(na3015_2), .IN4(1'b1), .IN5(na3017_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na4358_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y118     80'h00_0060_00_0000_0C06_FFA5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a230_4 ( .OUT(na230_2), .IN1(~na3017_2), .IN2(1'b0), .IN3(na3011_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x128y114     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a231_4 ( .OUT(na231_2), .IN1(na3017_2), .IN2(na3014_1), .IN3(~na3011_1), .IN4(~na4358_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x123y116     80'h00_0018_00_0000_0666_BC37
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(na220_2), .IN2(na3447_1), .IN3(1'b1), .IN4(na234_1), .IN5(1'b1), .IN6(~na3014_1), .IN7(~na236_1),
                     .IN8(na231_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y116     80'h00_0018_00_0040_0AD9_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_1 ( .OUT(na234_1), .IN1(1'b1), .IN2(na221_2), .IN3(~na222_2), .IN4(1'b1), .IN5(~na226_1), .IN6(1'b0), .IN7(na3449_2),
                     .IN8(~na230_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y113     80'h00_0018_00_0000_0C66_5A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_1 ( .OUT(na236_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3017_1), .IN6(1'b0), .IN7(~na3015_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x125y115     80'h00_0018_00_0000_0C88_39FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3016_1), .IN6(~na3014_1), .IN7(1'b0), .IN8(na4178_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y112     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_1 ( .OUT(na238_1), .IN1(~na220_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3017_2), .IN6(~na4357_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y114     80'h00_0018_00_0040_0AF8_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(1'b1), .IN2(na232_1), .IN3(1'b1), .IN4(~na1801_1), .IN5(na3451_1), .IN6(na1797_1), .IN7(na1799_1),
                     .IN8(~na4282_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y111     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a240_4 ( .OUT(na240_2), .IN1(~na220_2), .IN2(na221_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y112     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_1 ( .OUT(na241_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na242_2), .IN8(na231_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x134y111     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a242_4 ( .OUT(na242_2), .IN1(na3017_2), .IN2(na3013_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y109     80'h00_0018_00_0040_0A7E_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1), .IN1(1'b1), .IN2(na245_1), .IN3(1'b1), .IN4(~na4184_2), .IN5(na3452_2), .IN6(~na4187_2), .IN7(~na246_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y112     80'h00_0018_00_0040_0AF3_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a244_1 ( .OUT(na244_1), .IN1(1'b1), .IN2(~na1797_1), .IN3(~na1799_1), .IN4(1'b1), .IN5(~na4283_2), .IN6(~na232_1), .IN7(na3453_1),
                     .IN8(na1801_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y114     80'h00_0018_00_0040_0AF6_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a245_1 ( .OUT(na245_1), .IN1(1'b1), .IN2(~na1797_1), .IN3(1'b1), .IN4(~na1801_1), .IN5(na3454_2), .IN6(~na232_1), .IN7(~na1799_1),
                     .IN8(na4181_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x130y107     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_1 ( .OUT(na246_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3010_2), .IN6(~na247_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x131y112     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a247_4 ( .OUT(na247_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na236_1), .IN4(na227_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x128y110     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a248_1 ( .OUT(na248_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na222_2), .IN8(na230_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x115y110     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na252_1), .IN6(~na254_1), .IN7(na251_1), .IN8(na250_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y116     80'h00_0018_00_0040_0ADA_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a250_1 ( .OUT(na250_1), .IN1(na219_1), .IN2(1'b1), .IN3(~na236_1), .IN4(1'b1), .IN5(na226_1), .IN6(1'b1), .IN7(na3455_1),
                     .IN8(~na4184_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y109     80'h00_0018_00_0040_0AB5_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a251_1 ( .OUT(na251_1), .IN1(1'b1), .IN2(~na4182_2), .IN3(1'b1), .IN4(na4185_2), .IN5(~na220_2), .IN6(na3456_2), .IN7(1'b1),
                     .IN8(na4179_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y111     80'h00_0018_00_0040_0A7E_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1), .IN1(1'b1), .IN2(na245_1), .IN3(1'b1), .IN4(~na4184_2), .IN5(na3457_2), .IN6(~na253_2), .IN7(~na242_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x121y114     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a253_4 ( .OUT(na253_2), .IN1(na226_1), .IN2(1'b0), .IN3(na236_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y110     80'h00_0018_00_0040_0A79_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(na219_1), .IN2(1'b1), .IN3(1'b1), .IN4(na239_1), .IN5(~na220_2), .IN6(na3456_2), .IN7(na222_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x133y109     80'h00_0060_00_0000_0C06_FFE7
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a255_4 ( .OUT(na255_2), .IN1(na220_2), .IN2(na244_1), .IN3(~na222_2), .IN4(~na4185_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y112     80'h00_0018_00_0040_0A7A_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1), .IN1(na219_1), .IN2(1'b1), .IN3(1'b1), .IN4(na239_1), .IN5(na226_1), .IN6(~na253_2), .IN7(na236_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y110     80'h00_0018_00_0040_0A7E_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_1 ( .OUT(na258_1), .IN1(na219_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4186_2), .IN5(na3462_1), .IN6(~na244_1), .IN7(~na4355_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y111     80'h00_0018_00_0040_0A7E_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a259_1 ( .OUT(na259_1), .IN1(1'b1), .IN2(na245_1), .IN3(1'b1), .IN4(na239_1), .IN5(na3463_2), .IN6(~na4187_2), .IN7(~na240_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x116y81     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3465_1), .IN8(~na261_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y86     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a261_1 ( .OUT(na261_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4310_2), .IN5(~na3466_1), .IN6(1'b0), .IN7(~na3134_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x99y96     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a262_4 ( .OUT(na262_2), .IN1(~na2039_2), .IN2(~na16_2), .IN3(~na2007_2), .IN4(na19_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y108     80'h00_0018_00_0000_0666_066A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a263_1 ( .OUT(na263_1), .IN1(na252_1), .IN2(1'b0), .IN3(na259_1), .IN4(na258_1), .IN5(na264_1), .IN6(na254_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x115y107     80'h00_0018_00_0000_0666_A965
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a264_1 ( .OUT(na264_1), .IN1(~na267_1), .IN2(1'b0), .IN3(na268_1), .IN4(na250_1), .IN5(na217_1), .IN6(~na266_1), .IN7(na251_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y114     80'h00_0018_00_0040_0A71_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_1 ( .OUT(na266_1), .IN1(1'b1), .IN2(na4182_2), .IN3(1'b1), .IN4(na4185_2), .IN5(~na3452_2), .IN6(na4187_2), .IN7(na246_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y115     80'h00_0018_00_0040_0AE5_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(~na219_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4184_2), .IN5(1'b1), .IN6(na247_2), .IN7(~na240_2),
                     .IN8(na3470_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y113     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_1 ( .OUT(na268_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na255_2), .IN6(~na4188_2), .IN7(na4189_2), .IN8(na256_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y114     80'h00_0018_00_0040_0AD1_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_1 ( .OUT(na269_1), .IN1(1'b1), .IN2(na4182_2), .IN3(1'b1), .IN4(~na4176_2), .IN5(~na3463_2), .IN6(1'b0), .IN7(na240_2),
                     .IN8(na248_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y109     80'h00_0018_00_0040_0AE5_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a270_1 ( .OUT(na270_1), .IN1(1'b1), .IN2(~na245_1), .IN3(1'b1), .IN4(na4184_2), .IN5(1'b1), .IN6(na241_1), .IN7(~na246_1),
                     .IN8(na3472_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x118y84     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na273_1), .IN8(na3474_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y89     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na3475_2), .IN7(1'b0), .IN8(~na3135_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x114y93     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a274_4 ( .OUT(na274_2), .IN1(~na2040_1), .IN2(~na16_2), .IN3(~na2008_1), .IN4(na19_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x110y82     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a275_1 ( .OUT(na275_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na264_1), .IN6(1'b0), .IN7(na276_1), .IN8(na216_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y111     80'h00_0018_00_0000_0666_9996
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1), .IN1(na252_1), .IN2(na249_1), .IN3(na268_1), .IN4(~na258_1), .IN5(~na255_2), .IN6(na254_1), .IN7(na259_1),
                     .IN8(~na256_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x112y79     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3479_1), .IN8(~na279_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y80     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a279_1 ( .OUT(na279_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3480_2), .IN6(~na3136_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y92     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_1 ( .OUT(na280_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2041_2), .IN6(~na16_2), .IN7(~na2009_2),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y107     80'h00_0018_00_0000_0666_9963
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a281_1 ( .OUT(na281_1), .IN1(1'b0), .IN2(~na249_1), .IN3(na276_1), .IN4(na269_1), .IN5(na270_1), .IN6(~na284_1), .IN7(~na283_1),
                     .IN8(na216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y111     80'h00_0018_00_0040_0A74_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1), .IN1(1'b1), .IN2(~na244_1), .IN3(1'b1), .IN4(na4185_2), .IN5(na3483_2), .IN6(na253_2), .IN7(~na222_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y110     80'h00_0018_00_0040_0ADB_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(na219_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na239_1), .IN5(~na220_2), .IN6(1'b1), .IN7(na3484_1),
                     .IN8(~na4183_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x114y84     80'h00_0018_00_0000_0888_F33E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_1 ( .OUT(na285_1), .IN1(na21_2), .IN2(na3490_2), .IN3(1'b0), .IN4(~na286_1), .IN5(1'b0), .IN6(~na287_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y90     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a286_1 ( .OUT(na286_1), .IN1(1'b1), .IN2(na57_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na281_1), .IN8(na1978_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y92     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na288_1), .IN6(~na3486_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x103y97     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_1 ( .OUT(na288_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2042_1), .IN6(~na16_2), .IN7(~na2010_1),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y94     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a290_1 ( .OUT(na290_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2901_1), .IN6(na2362_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y94     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a292_1 ( .OUT(na292_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3137_1), .IN8(~na3492_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x106y79     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a293_1 ( .OUT(na293_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na276_1), .IN8(na4191_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y105     80'h00_0018_00_0000_0666_A999
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a294_1 ( .OUT(na294_1), .IN1(na267_1), .IN2(~na266_1), .IN3(~na283_1), .IN4(na269_1), .IN5(na270_1), .IN6(~na284_1), .IN7(na268_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x110y67     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a295_4 ( .OUT(na295_2), .IN1(~na21_2), .IN2(1'b0), .IN3(na3494_1), .IN4(~na296_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y78     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a296_1 ( .OUT(na296_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3495_2), .IN8(~na3138_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x102y84     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a297_4 ( .OUT(na297_2), .IN1(~na2043_2), .IN2(~na16_2), .IN3(~na2011_2), .IN4(na19_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y87     80'h00_0018_00_0000_0666_0695
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a298_1 ( .OUT(na298_1), .IN1(~na270_1), .IN2(1'b0), .IN3(na294_1), .IN4(~na269_1), .IN5(na217_1), .IN6(na249_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x109y68     80'h00_0018_00_0000_0888_F33E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a300_1 ( .OUT(na300_1), .IN1(na21_2), .IN2(na3503_1), .IN3(1'b0), .IN4(~na301_1), .IN5(1'b0), .IN6(~na302_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y76     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a301_1 ( .OUT(na301_1), .IN1(1'b1), .IN2(na57_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na298_1), .IN8(na1980_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y74     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a302_1 ( .OUT(na302_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3499_1), .IN6(~na303_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x103y74     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a303_4 ( .OUT(na303_2), .IN1(~na2044_1), .IN2(~na16_2), .IN3(~na2012_1), .IN4(na19_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y84     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a305_1 ( .OUT(na305_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2903_1), .IN8(na2364_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y78     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_1 ( .OUT(na307_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3505_2), .IN6(~na3139_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y93     80'h00_0018_00_0000_0666_A395
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a308_1 ( .OUT(na308_1), .IN1(~na267_1), .IN2(1'b0), .IN3(~na294_1), .IN4(na250_1), .IN5(1'b0), .IN6(~na266_1), .IN7(na251_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x114y79     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na310_1), .IN8(na3507_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y87     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a310_1 ( .OUT(na310_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3508_1), .IN6(~na3140_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x100y88     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2045_2), .IN6(~na16_2), .IN7(~na2013_2),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x109y79     80'h00_0018_00_0000_0666_6A09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_1 ( .OUT(na312_1), .IN1(~na264_1), .IN2(na249_1), .IN3(1'b0), .IN4(1'b0), .IN5(na217_1), .IN6(1'b0), .IN7(na294_1),
                     .IN8(na216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x108y71     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a313_4 ( .OUT(na313_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na314_1), .IN4(na3512_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a314_1 ( .OUT(na314_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3141_1), .IN6(~na3513_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x102y78     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a315_1 ( .OUT(na315_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2046_1), .IN6(~na16_2), .IN7(~na2014_1),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_1 ( .OUT(na316_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na324_1), .IN6(~na317_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x137y84     80'h00_0018_00_0000_0888_1545
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a317_1 ( .OUT(na317_1), .IN1(~na3519_1), .IN2(1'b1), .IN3(~na3516_1), .IN4(na3518_2), .IN5(~na3519_2), .IN6(1'b1), .IN7(~na320_1),
                     .IN8(~na319_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y90     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2994_2), .IN6(na2391_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y87     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_1 ( .OUT(na320_1), .IN1(1'b1), .IN2(na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na2930_2), .IN6(na1920_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y71     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(~na2416_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y77     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a323_4 ( .OUT(na323_2), .IN1(~na21_2), .IN2(na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x103y95     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1), .IN1(na21_2), .IN2(~na2095_2), .IN3(na26_2), .IN4(~na1967_2), .IN5(~na2031_2), .IN6(~na16_2), .IN7(~na1999_2),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y77     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na328_1), .IN8(~na3523_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x118y93     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1), .IN1(na21_2), .IN2(~na2096_1), .IN3(~na2000_1), .IN4(na19_1), .IN5(~na2032_1), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na1968_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x125y86     80'h00_0018_00_0000_0CEE_A300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a332_1 ( .OUT(na332_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na16_2), .IN7(na3529_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y93     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a334_1 ( .OUT(na334_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2392_2), .IN8(na2995_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y89     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na1921_2), .IN6(na2931_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y78     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a336_1 ( .OUT(na336_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3531_1), .IN8(~na339_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x110y94     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a339_1 ( .OUT(na339_1), .IN1(na21_2), .IN2(~na2097_2), .IN3(~na2001_2), .IN4(na19_1), .IN5(~na2033_2), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na1969_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y85     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2393_1), .IN8(na2996_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y84     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a344_1 ( .OUT(na344_1), .IN1(1'b1), .IN2(na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na2932_2), .IN6(na1922_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a345_1 ( .OUT(na345_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na348_1), .IN6(~na3540_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x105y95     80'h00_0018_00_0000_0888_7BDB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_1 ( .OUT(na348_1), .IN1(na4168_2), .IN2(~na1970_1), .IN3(~na2002_1), .IN4(na19_1), .IN5(na21_2), .IN6(~na2098_1), .IN7(~na4163_2),
                     .IN8(~na2034_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y88     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2997_1), .IN6(na2394_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y85     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2933_1), .IN8(na1923_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y76     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4172_2), .IN5(1'b0), .IN6(~na355_1), .IN7(1'b0), .IN8(~na360_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x137y68     80'h00_0018_00_0000_0888_511C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1), .IN1(1'b1), .IN2(na3550_2), .IN3(~na3551_1), .IN4(~na3548_2), .IN5(~na357_1), .IN6(~na358_1), .IN7(~na3551_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y79     80'h00_0018_00_0040_0A50_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b1), .IN2(na4164_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(na2998_2), .IN6(1'b0), .IN7(na2395_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y78     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b1), .IN2(na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na2934_2), .IN6(na1924_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y86     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a360_1 ( .OUT(na360_1), .IN1(na21_2), .IN2(~na2099_2), .IN3(na26_2), .IN4(~na1971_2), .IN5(~na2035_2), .IN6(~na16_2), .IN7(~na2003_2),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y74     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3555_1), .IN8(~na366_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x104y76     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1), .IN1(na21_2), .IN2(~na2100_1), .IN3(~na2004_1), .IN4(na19_1), .IN5(~na2036_1), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na1972_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y77     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_1 ( .OUT(na370_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2396_2), .IN6(na2999_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y74     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a371_1 ( .OUT(na371_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2935_1), .IN8(na1925_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y76     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a372_1 ( .OUT(na372_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na373_1), .IN8(~na378_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y75     80'h00_0018_00_0000_0888_5145
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a373_1 ( .OUT(na373_1), .IN1(~na3566_1), .IN2(1'b1), .IN3(~na3563_1), .IN4(na3565_1), .IN5(~na3566_2), .IN6(~na375_1), .IN7(~na376_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y84     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_1 ( .OUT(na375_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3000_2), .IN8(na2397_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y83     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a376_1 ( .OUT(na376_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na1926_1), .IN6(na2936_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x108y84     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(na21_2), .IN2(~na2101_2), .IN3(~na2005_2), .IN4(na19_1), .IN5(~na2037_2), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na1973_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y77     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4172_2), .IN5(~na382_1), .IN6(1'b0), .IN7(~na387_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x131y69     80'h00_0018_00_0000_0888_5345
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_1 ( .OUT(na382_1), .IN1(~na4397_2), .IN2(1'b1), .IN3(~na3570_1), .IN4(na386_2), .IN5(1'b1), .IN6(~na385_1), .IN7(~na384_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y79     80'h00_0018_00_0040_0AA0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a384_1 ( .OUT(na384_1), .IN1(1'b1), .IN2(~na4164_2), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(na2398_2), .IN7(1'b0),
                     .IN8(na3001_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y78     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a385_1 ( .OUT(na385_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2937_1), .IN8(na1927_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x126y74     80'h00_0060_00_0000_0C0E_FF0B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a386_4 ( .OUT(na386_2), .IN1(na3572_1), .IN2(~na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x102y75     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a387_1 ( .OUT(na387_1), .IN1(na21_2), .IN2(~na2102_1), .IN3(na26_2), .IN4(~na1974_1), .IN5(~na2038_1), .IN6(~na16_2), .IN7(~na2006_1),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y79     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a390_1 ( .OUT(na390_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3576_1), .IN6(~na391_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x137y88     80'h00_0018_00_0000_0888_3123
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1), .IN1(1'b1), .IN2(~na3580_1), .IN3(na3579_1), .IN4(~na3577_2), .IN5(~na393_1), .IN6(~na3580_2), .IN7(1'b1),
                     .IN8(~na394_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y93     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2922_2), .IN8(na3066_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y88     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a394_1 ( .OUT(na394_1), .IN1(1'b1), .IN2(na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na2335_1), .IN6(na3082_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y79     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a398_1 ( .OUT(na398_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4172_2), .IN5(1'b0), .IN6(~na404_1), .IN7(1'b0), .IN8(~na399_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y90     80'h00_0018_00_0000_0888_1A53
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b1), .IN2(~na402_1), .IN3(~na3585_1), .IN4(1'b1), .IN5(na403_1), .IN6(1'b1), .IN7(~na3585_2),
                     .IN8(~na401_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y94     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a401_1 ( .OUT(na401_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2923_1), .IN6(na3067_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y88     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a402_1 ( .OUT(na402_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3083_2), .IN8(na2336_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y91     80'h00_0018_00_0040_0A5F_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(~na2344_2), .IN6(1'b1), .IN7(~na3043_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x117y96     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a404_1 ( .OUT(na404_1), .IN1(na21_2), .IN2(~na2056_1), .IN3(~na1992_1), .IN4(na19_1), .IN5(~na2024_1), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na1960_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y77     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a407_1 ( .OUT(na407_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na408_1), .IN8(~na413_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x136y71     80'h00_0018_00_0000_0888_5123
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1), .IN1(1'b1), .IN2(~na3593_1), .IN3(na3592_1), .IN4(~na3590_2), .IN5(~na411_1), .IN6(~na3593_2), .IN7(~na410_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y83     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a410_1 ( .OUT(na410_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3068_2), .IN8(na2924_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y79     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3084_2), .IN8(na2337_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x110y92     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1), .IN1(na21_2), .IN2(~na2057_2), .IN3(~na1993_2), .IN4(na19_1), .IN5(~na2025_2), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na1961_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y77     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na417_1), .IN6(~na422_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x135y81     80'h00_0018_00_0000_0888_1233
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1), .IN1(1'b1), .IN2(~na3597_2), .IN3(1'b1), .IN4(~na3599_2), .IN5(na3598_1), .IN6(~na420_1), .IN7(~na421_1),
                     .IN8(~na3599_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y88     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a420_1 ( .OUT(na420_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2925_1), .IN6(na3069_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y85     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3085_1), .IN8(na2338_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y94     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a422_1 ( .OUT(na422_1), .IN1(na21_2), .IN2(~na2058_1), .IN3(na26_2), .IN4(~na1962_1), .IN5(~na2026_1), .IN6(~na16_2), .IN7(~na1994_1),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y74     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na431_1), .IN6(~na426_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y66     80'h00_0018_00_0000_0888_3154
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a426_1 ( .OUT(na426_1), .IN1(~na3607_2), .IN2(na3606_1), .IN3(~na3604_2), .IN4(1'b1), .IN5(~na3607_1), .IN6(~na429_1), .IN7(1'b1),
                     .IN8(~na428_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y78     80'h00_0018_00_0040_0A50_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a428_1 ( .OUT(na428_1), .IN1(1'b1), .IN2(na4164_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(na3070_2), .IN6(1'b0), .IN7(na2926_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y74     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na3086_2), .IN6(na2339_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y85     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1), .IN1(na21_2), .IN2(~na2059_2), .IN3(na26_2), .IN4(~na1963_2), .IN5(~na2027_2), .IN6(~na16_2), .IN7(~na1995_2),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y73     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a434_1 ( .OUT(na434_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3611_1), .IN8(~na435_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y66     80'h00_0018_00_0000_0888_5123
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1), .IN1(1'b1), .IN2(~na3615_1), .IN3(na3614_2), .IN4(~na3612_1), .IN5(~na438_1), .IN6(~na3615_2), .IN7(~na437_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y75     80'h00_0018_00_0040_0AA0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1), .IN1(1'b1), .IN2(~na4164_2), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(na2927_1), .IN7(1'b0),
                     .IN8(na3071_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y71     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na3087_1), .IN6(na2340_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y75     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na448_1), .IN6(~na443_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y68     80'h00_0018_00_0000_0888_2513
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1), .IN1(1'b1), .IN2(~na3620_1), .IN3(~na446_1), .IN4(~na3622_2), .IN5(~na447_1), .IN6(1'b1), .IN7(na3621_2),
                     .IN8(~na3622_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y79     80'h00_0018_00_0040_0AA0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a446_1 ( .OUT(na446_1), .IN1(1'b1), .IN2(~na4164_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(na3072_2), .IN7(1'b0),
                     .IN8(na2928_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y75     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a447_1 ( .OUT(na447_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na3088_2), .IN6(na2341_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y83     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a448_1 ( .OUT(na448_1), .IN1(na21_2), .IN2(~na2061_2), .IN3(~na1997_2), .IN4(na19_1), .IN5(~na2029_2), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na1965_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y73     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4172_2), .IN5(~na457_1), .IN6(1'b0), .IN7(~na452_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x130y67     80'h00_0018_00_0000_0888_15F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(~na3627_2), .IN2(na456_1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3627_1), .IN6(1'b1), .IN7(~na454_1),
                     .IN8(~na455_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y75     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a454_1 ( .OUT(na454_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2929_1), .IN8(na3073_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y74     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na3089_1), .IN6(na2342_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x127y72     80'h00_0018_00_0000_0CEE_0B00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a456_1 ( .OUT(na456_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3629_1), .IN6(~na16_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x103y73     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_1 ( .OUT(na457_1), .IN1(na21_2), .IN2(~na2062_1), .IN3(na26_2), .IN4(~na1966_1), .IN5(~na2030_1), .IN6(~na16_2), .IN7(~na1998_1),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y80     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a460_1 ( .OUT(na460_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na463_1), .IN6(~na3633_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y95     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a463_1 ( .OUT(na463_1), .IN1(na21_2), .IN2(~na2047_2), .IN3(~na1983_2), .IN4(na19_1), .IN5(~na2015_2), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na3186_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y93     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2938_2), .IN6(na2327_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y90     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a468_1 ( .OUT(na468_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na3074_2), .IN6(na2367_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y80     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a469_1 ( .OUT(na469_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3641_1), .IN6(~na470_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y92     80'h00_0018_00_0000_0888_141F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na3642_1), .IN4(~na3644_2), .IN5(~na473_1), .IN6(na3643_2), .IN7(~na474_1),
                     .IN8(~na3644_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y95     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a473_1 ( .OUT(na473_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2939_1), .IN6(na2328_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y91     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a474_1 ( .OUT(na474_1), .IN1(1'b1), .IN2(na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na2368_2), .IN6(na3075_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y80     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na480_1), .IN6(~na3650_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x111y93     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a480_1 ( .OUT(na480_1), .IN1(na21_2), .IN2(~na2049_2), .IN3(~na1985_2), .IN4(na19_1), .IN5(~na2017_2), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na3188_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y87     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_1 ( .OUT(na484_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2329_1), .IN8(na2940_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y84     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a485_1 ( .OUT(na485_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na3076_2), .IN6(na2369_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y77     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na487_1), .IN8(~na3659_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y93     80'h00_0018_00_0000_0888_7BDB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a487_1 ( .OUT(na487_1), .IN1(na4168_2), .IN2(~na3189_1), .IN3(~na1986_1), .IN4(na19_1), .IN5(na21_2), .IN6(~na2050_1), .IN7(~na4163_2),
                     .IN8(~na2018_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y87     80'h00_0018_00_0040_0A3F_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(~na3061_1), .IN6(~na2378_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y92     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_1 ( .OUT(na493_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2941_1), .IN6(na2330_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y86     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a494_1 ( .OUT(na494_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2370_2), .IN8(na3077_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y75     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na496_1), .IN6(~na501_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x135y71     80'h00_0018_00_0000_0888_5154
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a496_1 ( .OUT(na496_1), .IN1(~na3668_1), .IN2(na3667_2), .IN3(~na3665_1), .IN4(1'b1), .IN5(~na3668_2), .IN6(~na499_1), .IN7(~na498_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y81     80'h00_0018_00_0040_0A50_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a498_1 ( .OUT(na498_1), .IN1(1'b1), .IN2(na4164_2), .IN3(1'b1), .IN4(na4310_2), .IN5(na2331_1), .IN6(1'b0), .IN7(na2942_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y80     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a499_1 ( .OUT(na499_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(na26_2), .IN4(1'b1), .IN5(na3078_2), .IN6(na2371_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y86     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1), .IN1(na21_2), .IN2(~na2051_2), .IN3(na26_2), .IN4(~na3190_2), .IN5(~na2019_2), .IN6(~na16_2), .IN7(~na1987_2),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y75     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a504_1 ( .OUT(na504_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4172_2), .IN5(1'b0), .IN6(~na510_1), .IN7(1'b0), .IN8(~na3672_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y80     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a508_1 ( .OUT(na508_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2943_1), .IN6(na2332_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y76     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a509_1 ( .OUT(na509_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2372_2), .IN8(na3079_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x105y78     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a510_1 ( .OUT(na510_1), .IN1(na21_2), .IN2(~na2052_1), .IN3(~na1988_1), .IN4(na19_1), .IN5(~na2020_1), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na3191_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y75     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a513_1 ( .OUT(na513_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4172_2), .IN5(1'b0), .IN6(~na516_1), .IN7(1'b0), .IN8(~na3680_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y84     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a516_1 ( .OUT(na516_1), .IN1(na21_2), .IN2(~na2053_2), .IN3(~na1989_2), .IN4(na19_1), .IN5(~na2021_2), .IN6(~na16_2), .IN7(na26_2),
                     .IN8(~na3192_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y90     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a520_1 ( .OUT(na520_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2944_2), .IN6(na2333_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y86     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a521_1 ( .OUT(na521_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2373_1), .IN8(na3080_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y69     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a522_1 ( .OUT(na522_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na523_1), .IN8(~na528_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y79     80'h00_0018_00_0000_0888_C155
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1), .IN1(~na3689_1), .IN2(1'b1), .IN3(~na526_1), .IN4(1'b1), .IN5(~na3689_2), .IN6(~na525_1), .IN7(1'b1),
                     .IN8(na527_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y88     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(na2945_1), .IN6(na2334_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y83     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a526_1 ( .OUT(na526_1), .IN1(1'b1), .IN2(na2416_2), .IN3(~na26_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2374_2), .IN8(na3081_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y82     80'h00_0018_00_0040_0A3F_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a527_1 ( .OUT(na527_1), .IN1(1'b1), .IN2(na2416_2), .IN3(na4165_2), .IN4(1'b1), .IN5(~na2382_2), .IN6(~na3065_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x104y78     80'h00_0018_00_0000_0888_D7BB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a528_1 ( .OUT(na528_1), .IN1(na21_2), .IN2(~na2054_1), .IN3(na26_2), .IN4(~na3193_1), .IN5(~na2022_1), .IN6(~na16_2), .IN7(~na1990_1),
                     .IN8(na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y69     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a531_4 ( .OUT(na531_2), .IN1(na532_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na536_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y67     80'h00_0018_00_0040_0A37_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a532_1 ( .OUT(na532_1), .IN1(1'b1), .IN2(~na1957_2), .IN3(na1958_1), .IN4(1'b1), .IN5(~na533_1), .IN6(~na534_2), .IN7(1'b1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x131y67     80'h00_0018_00_0040_0CFA_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1), .IN1(1'b1), .IN2(~na3694_2), .IN3(1'b1), .IN4(~na3150_2), .IN5(~na4381_2), .IN6(1'b1), .IN7(na3151_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y102     80'h00_0060_00_0000_0C08_FFC8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a534_4 ( .OUT(na534_2), .IN1(na4299_2), .IN2(na535_2), .IN3(1'b1), .IN4(na1938_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y98     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a535_4 ( .OUT(na535_2), .IN1(~na1935_1), .IN2(~na1937_2), .IN3(~na4298_2), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y70     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a536_4 ( .OUT(na536_2), .IN1(~na537_1), .IN2(1'b1), .IN3(na1958_1), .IN4(~na3695_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y71     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a537_1 ( .OUT(na537_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4296_2), .IN6(~na1929_1), .IN7(na538_1),
                     .IN8(na1932_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y77     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a538_1 ( .OUT(na538_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1930_1), .IN8(~na1932_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y80     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a539_4 ( .OUT(na539_2), .IN1(1'b1), .IN2(~na4392_2), .IN3(~na3223_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x141y70     80'h00_0018_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a540_1 ( .OUT(na540_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1958_1), .IN4(1'b1), .IN5(1'b0), .IN6(na3696_1), .IN7(1'b0), .IN8(~na541_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y70     80'h00_0018_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a541_1 ( .OUT(na541_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na537_1), .IN6(na1957_2), .IN7(1'b1), .IN8(~na3695_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y104     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a542_1 ( .OUT(na542_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2578_2), .IN6(na2191_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x107y92     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a543_4 ( .OUT(na543_2), .IN1(1'b0), .IN2(~na3285_2), .IN3(~na3151_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y103     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a544_1 ( .OUT(na544_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2192_1), .IN6(na2579_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y91     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a545_1 ( .OUT(na545_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2580_2), .IN6(na2193_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y108     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a546_1 ( .OUT(na546_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2581_1), .IN6(na2194_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y86     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a547_1 ( .OUT(na547_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2195_2), .IN6(na2582_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y90     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a548_1 ( .OUT(na548_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2583_1), .IN6(na2196_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y87     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a549_1 ( .OUT(na549_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2584_2), .IN6(na2197_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y75     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a550_1 ( .OUT(na550_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2585_1), .IN6(na2198_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y112     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a551_1 ( .OUT(na551_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2586_2), .IN6(na2199_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y104     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a552_1 ( .OUT(na552_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2200_1), .IN6(na2587_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y108     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a553_1 ( .OUT(na553_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2588_2), .IN8(na2201_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y111     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a554_1 ( .OUT(na554_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2589_1), .IN6(na2202_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y96     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a555_1 ( .OUT(na555_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2590_2), .IN6(na2203_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y71     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a556_1 ( .OUT(na556_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2204_1), .IN6(na2591_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y100     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a557_1 ( .OUT(na557_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2592_2), .IN6(na2205_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y70     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a558_1 ( .OUT(na558_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2593_1), .IN6(na2206_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y109     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a559_1 ( .OUT(na559_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2594_1), .IN6(na2207_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y101     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a560_1 ( .OUT(na560_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2595_1), .IN8(na2208_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y97     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a561_1 ( .OUT(na561_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2596_2), .IN6(na2209_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y110     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a562_1 ( .OUT(na562_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2597_1), .IN6(na2210_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y93     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a563_1 ( .OUT(na563_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2598_2), .IN8(na2211_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y70     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a564_1 ( .OUT(na564_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2212_2), .IN6(na2599_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y85     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a565_1 ( .OUT(na565_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2213_1), .IN8(na2600_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y84     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a566_1 ( .OUT(na566_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2601_1), .IN6(na2214_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y109     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2159_2), .IN8(na2602_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y104     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a568_1 ( .OUT(na568_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2603_1), .IN6(na2160_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y107     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_1 ( .OUT(na569_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2604_2), .IN6(na2161_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y109     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a570_1 ( .OUT(na570_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2605_1), .IN8(na2162_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y105     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a571_1 ( .OUT(na571_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2606_2), .IN8(na2163_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y90     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a572_1 ( .OUT(na572_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2607_1), .IN8(na2164_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y97     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a573_1 ( .OUT(na573_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2608_2), .IN6(na2165_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y89     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a574_1 ( .OUT(na574_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2609_1), .IN8(na2166_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y108     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a575_1 ( .OUT(na575_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3194_2), .IN6(na2730_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y103     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a576_1 ( .OUT(na576_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2731_1), .IN6(na3195_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y103     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_1 ( .OUT(na577_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3196_2), .IN6(na2732_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y111     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a578_1 ( .OUT(na578_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2733_1), .IN8(na3197_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y99     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_1 ( .OUT(na579_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3198_2), .IN6(na2734_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y87     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a580_1 ( .OUT(na580_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2735_1), .IN6(na3199_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y99     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_1 ( .OUT(na581_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3200_2), .IN6(na2736_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y92     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a582_1 ( .OUT(na582_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2737_1), .IN8(na3201_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y108     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_1 ( .OUT(na583_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3142_1), .IN6(na2706_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y104     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a584_1 ( .OUT(na584_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3143_1), .IN6(na2707_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x108y93     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_1 ( .OUT(na585_1), .IN1(na3144_2), .IN2(na2708_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y107     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a586_1 ( .OUT(na586_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2709_1), .IN8(na3145_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x96y90     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_1 ( .OUT(na587_1), .IN1(na2710_2), .IN2(na3146_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x99y82     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a588_1 ( .OUT(na588_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2711_2), .IN8(na3147_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x97y96     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a589_1 ( .OUT(na589_1), .IN1(na2712_2), .IN2(na3148_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y74     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a590_1 ( .OUT(na590_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2713_1), .IN6(na3149_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x105y111     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a591_1 ( .OUT(na591_1), .IN1(na2714_2), .IN2(na1912_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y104     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a592_1 ( .OUT(na592_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2715_1), .IN6(na1913_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y109     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a593_1 ( .OUT(na593_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1914_1), .IN6(na2716_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y112     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_1 ( .OUT(na594_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2717_1), .IN6(na1915_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y98     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a595_1 ( .OUT(na595_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1916_1), .IN6(na2718_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x104y71     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a596_1 ( .OUT(na596_1), .IN1(na1917_2), .IN2(na2719_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y93     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a597_1 ( .OUT(na597_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2720_2), .IN6(na1918_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y78     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a598_1 ( .OUT(na598_1), .IN1(na2721_1), .IN2(na1919_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y108     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a599_1 ( .OUT(na599_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2722_2), .IN6(na1903_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y99     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a600_1 ( .OUT(na600_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2723_1), .IN8(na1904_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y104     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a601_1 ( .OUT(na601_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2724_2), .IN8(na1905_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y110     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a602_1 ( .OUT(na602_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1906_1), .IN6(na2725_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x101y101     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a603_1 ( .OUT(na603_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2726_2), .IN4(na1907_2), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y76     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a604_1 ( .OUT(na604_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2727_1), .IN6(na1908_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x111y89     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a605_1 ( .OUT(na605_1), .IN1(na2728_2), .IN2(na1909_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y84     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a606_1 ( .OUT(na606_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1910_1), .IN6(na2729_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y103     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a607_1 ( .OUT(na607_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2482_2), .IN8(na2071_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y103     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a608_1 ( .OUT(na608_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2072_1), .IN6(na2483_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y82     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a609_1 ( .OUT(na609_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2484_2), .IN8(na2073_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y107     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a610_1 ( .OUT(na610_1), .IN1(na2074_1), .IN2(na2485_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y86     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a611_1 ( .OUT(na611_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2486_2), .IN8(na2075_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y83     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a612_1 ( .OUT(na612_1), .IN1(na2487_1), .IN2(na2076_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y89     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a613_1 ( .OUT(na613_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2077_2), .IN8(na2488_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y71     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a614_1 ( .OUT(na614_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2078_1), .IN6(na2489_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y112     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a615_1 ( .OUT(na615_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2490_2), .IN8(na2079_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y101     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a616_1 ( .OUT(na616_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2491_1), .IN8(na2080_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x120y111     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a617_1 ( .OUT(na617_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2081_2), .IN4(na2492_2), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y106     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a618_1 ( .OUT(na618_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2493_1), .IN6(na2082_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x114y91     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a619_1 ( .OUT(na619_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2083_2), .IN4(na2494_2), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y80     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a620_1 ( .OUT(na620_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2495_1), .IN8(na2084_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y99     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a621_1 ( .OUT(na621_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2085_2), .IN8(na2496_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y75     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a622_1 ( .OUT(na622_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2497_1), .IN8(na2086_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y106     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a623_1 ( .OUT(na623_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1949_2), .IN8(na2498_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x125y101     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a624_1 ( .OUT(na624_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1950_1), .IN4(na2499_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y102     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a625_1 ( .OUT(na625_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1951_2), .IN6(na2500_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x112y107     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a626_1 ( .OUT(na626_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2501_1), .IN4(na1952_1), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y85     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a627_1 ( .OUT(na627_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1953_2), .IN6(na2502_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y69     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a628_1 ( .OUT(na628_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2503_1), .IN8(na1954_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y88     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a629_1 ( .OUT(na629_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1955_2), .IN6(na2504_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y83     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a630_1 ( .OUT(na630_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2505_2), .IN8(na1956_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y107     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a631_1 ( .OUT(na631_1), .IN1(na3225_1), .IN2(na2506_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y110     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a632_1 ( .OUT(na632_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3226_2), .IN8(na2507_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x106y107     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a633_1 ( .OUT(na633_1), .IN1(na3227_1), .IN2(na2508_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y103     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a634_1 ( .OUT(na634_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2509_1), .IN8(na3228_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y101     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2510_2), .IN6(na3229_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y97     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a636_1 ( .OUT(na636_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2511_1), .IN6(na3230_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y106     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a637_1 ( .OUT(na637_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2512_2), .IN6(na3231_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y96     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a638_1 ( .OUT(na638_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3232_2), .IN4(na2513_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y107     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_1 ( .OUT(na639_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2143_2), .IN6(na2514_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x101y107     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a640_1 ( .OUT(na640_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2515_1), .IN4(na2144_1), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y87     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_1 ( .OUT(na641_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2516_2), .IN6(na2145_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y114     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a642_1 ( .OUT(na642_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2517_1), .IN6(na2146_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y87     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a643_1 ( .OUT(na643_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2147_2), .IN8(na2518_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x99y85     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a644_1 ( .OUT(na644_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2519_1), .IN6(na2148_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y87     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a645_1 ( .OUT(na645_1), .IN1(na2149_2), .IN2(na2520_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y74     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a646_1 ( .OUT(na646_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2150_1), .IN6(na2521_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x108y113     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a647_1 ( .OUT(na647_1), .IN1(na2522_2), .IN2(na2151_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y104     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a648_1 ( .OUT(na648_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2523_1), .IN6(na2152_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y106     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a649_1 ( .OUT(na649_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2524_2), .IN8(na2153_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y112     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a650_1 ( .OUT(na650_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2525_1), .IN6(na2154_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y96     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a651_1 ( .OUT(na651_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2526_2), .IN8(na2155_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x98y71     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a652_1 ( .OUT(na652_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2156_1), .IN4(na2527_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y104     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a653_1 ( .OUT(na653_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2157_2), .IN6(na2528_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x92y80     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a654_1 ( .OUT(na654_1), .IN1(na2529_1), .IN2(na2158_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y114     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2530_2), .IN6(na2103_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y100     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a656_1 ( .OUT(na656_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2104_1), .IN6(na2531_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y110     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a657_1 ( .OUT(na657_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2105_2), .IN6(na2532_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y114     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a658_1 ( .OUT(na658_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2533_1), .IN6(na2106_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x112y91     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a659_1 ( .OUT(na659_1), .IN1(na2107_2), .IN2(na2534_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y73     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a660_1 ( .OUT(na660_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2535_2), .IN6(na2108_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x115y86     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a661_1 ( .OUT(na661_1), .IN1(na2536_2), .IN2(na2109_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y85     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a662_1 ( .OUT(na662_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2110_1), .IN6(na2537_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y111     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a663_1 ( .OUT(na663_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2538_2), .IN6(na2063_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y104     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a664_1 ( .OUT(na664_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2539_1), .IN8(na2064_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y114     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a665_1 ( .OUT(na665_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2065_2), .IN8(na2540_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x98y112     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a666_1 ( .OUT(na666_1), .IN1(na2066_1), .IN2(na2541_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y106     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a667_1 ( .OUT(na667_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2542_2), .IN8(na2067_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y94     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a668_1 ( .OUT(na668_1), .IN1(na2543_1), .IN2(na2068_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y102     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a669_1 ( .OUT(na669_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2544_2), .IN8(na2069_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y93     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a670_1 ( .OUT(na670_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2070_1), .IN6(na2545_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y106     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a671_1 ( .OUT(na671_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2546_2), .IN6(na2111_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y104     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a672_1 ( .OUT(na672_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2112_1), .IN6(na2547_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x96y84     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a673_1 ( .OUT(na673_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2113_2), .IN4(na2548_2), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y112     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a674_1 ( .OUT(na674_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2549_1), .IN6(na2114_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y84     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a675_1 ( .OUT(na675_1), .IN1(na2115_2), .IN2(na2550_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y85     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a676_1 ( .OUT(na676_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2551_1), .IN8(na2116_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y86     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a677_1 ( .OUT(na677_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2552_2), .IN6(na2117_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a678_1 ( .OUT(na678_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2553_1), .IN6(na2118_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y114     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a679_1 ( .OUT(na679_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2119_2), .IN6(na2554_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x138y108     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a680_1 ( .OUT(na680_1), .IN1(na2120_1), .IN2(na2555_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y101     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a681_1 ( .OUT(na681_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2121_2), .IN6(na2556_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x101y114     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a682_1 ( .OUT(na682_1), .IN1(na2557_1), .IN2(na2122_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y96     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a683_1 ( .OUT(na683_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2558_2), .IN8(na2123_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y78     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a684_1 ( .OUT(na684_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2559_1), .IN6(na2124_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y102     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2560_2), .IN6(na2125_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y78     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a686_1 ( .OUT(na686_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2561_1), .IN8(na2126_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x121y108     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a687_1 ( .OUT(na687_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2562_2), .IN4(na2127_2), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y100     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a688_1 ( .OUT(na688_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2563_1), .IN6(na2128_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x110y109     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a689_1 ( .OUT(na689_1), .IN1(na2564_1), .IN2(na2129_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y112     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a690_1 ( .OUT(na690_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2130_1), .IN8(na2565_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y90     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a691_1 ( .OUT(na691_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2566_2), .IN6(na2131_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y69     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a692_1 ( .OUT(na692_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2567_1), .IN6(na2132_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y83     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a693_1 ( .OUT(na693_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2568_2), .IN6(na2133_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y86     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a694_1 ( .OUT(na694_1), .IN1(na2569_1), .IN2(na2134_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y112     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2570_2), .IN6(na2135_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x120y106     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a696_1 ( .OUT(na696_1), .IN1(na2136_2), .IN2(na2571_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y113     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a697_1 ( .OUT(na697_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2572_2), .IN6(na2137_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y113     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a698_1 ( .OUT(na698_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2573_1), .IN6(na2138_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y106     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a699_1 ( .OUT(na699_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2139_2), .IN6(na2574_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y93     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a700_1 ( .OUT(na700_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2575_1), .IN6(na2140_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y99     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a701_1 ( .OUT(na701_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2141_2), .IN4(na2576_2), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y94     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2142_1), .IN6(na2577_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y105     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1), .IN1(na2610_2), .IN2(na2215_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y105     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a704_1 ( .OUT(na704_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2216_2), .IN6(na2611_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y89     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a705_1 ( .OUT(na705_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2612_2), .IN8(na2217_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y109     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a706_1 ( .OUT(na706_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2218_2), .IN6(na2613_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y92     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2614_2), .IN6(na2219_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x93y77     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a708_1 ( .OUT(na708_1), .IN1(na2615_1), .IN2(na2220_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y94     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2616_2), .IN6(na2221_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x96y71     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a710_1 ( .OUT(na710_1), .IN1(na2617_1), .IN2(na2222_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y112     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2618_2), .IN8(na2167_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y104     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a712_1 ( .OUT(na712_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2619_1), .IN6(na2168_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y107     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a713_1 ( .OUT(na713_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2620_2), .IN8(na2169_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y104     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a714_1 ( .OUT(na714_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2621_1), .IN8(na2170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x121y91     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a715_1 ( .OUT(na715_1), .IN1(na2171_2), .IN2(na2622_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y70     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a716_1 ( .OUT(na716_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2623_2), .IN6(na2172_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x107y103     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a717_1 ( .OUT(na717_1), .IN1(na2173_2), .IN2(na2624_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y70     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a718_1 ( .OUT(na718_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2625_1), .IN8(na2174_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y108     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2626_2), .IN6(na2175_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y100     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a720_1 ( .OUT(na720_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2627_1), .IN6(na2176_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y105     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2628_2), .IN6(na2177_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x114y99     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a722_1 ( .OUT(na722_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2178_1), .IN4(na2629_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y86     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2630_2), .IN6(na2179_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x106y70     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a724_1 ( .OUT(na724_1), .IN1(na2631_1), .IN2(na2180_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y92     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a725_1 ( .OUT(na725_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2181_2), .IN6(na2632_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y86     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a726_1 ( .OUT(na726_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2182_1), .IN8(na2633_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y105     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2183_2), .IN6(na2634_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y103     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a728_1 ( .OUT(na728_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2635_1), .IN8(na2184_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x103y109     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a729_1 ( .OUT(na729_1), .IN1(na2185_2), .IN2(na2636_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y114     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a730_1 ( .OUT(na730_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2637_1), .IN6(na2186_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y104     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1), .IN1(na2187_2), .IN2(na2638_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y85     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a732_1 ( .OUT(na732_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2639_1), .IN8(na2188_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y100     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a733_1 ( .OUT(na733_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2640_2), .IN6(na2189_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y87     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a734_1 ( .OUT(na734_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2641_1), .IN6(na2190_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y108     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a735_1 ( .OUT(na735_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2642_2), .IN6(na2239_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x110y106     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a736_1 ( .OUT(na736_1), .IN1(na2643_1), .IN2(na2240_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y89     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2644_2), .IN6(na2241_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x92y113     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a738_1 ( .OUT(na738_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2645_1), .IN4(na2242_2), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y92     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2243_1), .IN6(na2646_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y82     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a740_1 ( .OUT(na740_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2647_1), .IN6(na2244_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y97     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a741_1 ( .OUT(na741_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2245_1), .IN6(na2648_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y69     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a742_1 ( .OUT(na742_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2246_2), .IN6(na2649_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x105y113     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a743_1 ( .OUT(na743_1), .IN1(na2247_1), .IN2(na2650_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y106     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a744_1 ( .OUT(na744_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2248_2), .IN8(na2651_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x117y112     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a745_1 ( .OUT(na745_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2249_1), .IN4(na2652_2), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y112     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a746_1 ( .OUT(na746_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2653_2), .IN6(na2250_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y105     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a747_1 ( .OUT(na747_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2654_2), .IN6(na2251_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y70     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a748_1 ( .OUT(na748_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2655_1), .IN6(na2252_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y100     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a749_1 ( .OUT(na749_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2656_2), .IN8(na2253_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x92y75     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a750_1 ( .OUT(na750_1), .IN1(na2657_1), .IN2(na2254_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y108     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a751_1 ( .OUT(na751_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2658_2), .IN8(na2255_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x130y102     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a752_1 ( .OUT(na752_1), .IN1(na2256_2), .IN2(na2659_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y110     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_1 ( .OUT(na753_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2660_2), .IN6(na2257_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y111     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a754_1 ( .OUT(na754_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2661_1), .IN6(na2258_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y89     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a755_1 ( .OUT(na755_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2662_2), .IN6(na2259_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y68     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a756_1 ( .OUT(na756_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2260_2), .IN6(na2663_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x111y88     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a757_1 ( .OUT(na757_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2664_2), .IN4(na2261_1), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y81     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a758_1 ( .OUT(na758_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2665_1), .IN6(na2262_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x95y113     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_1 ( .OUT(na759_1), .IN1(na2263_1), .IN2(na2666_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y106     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a760_1 ( .OUT(na760_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2667_1), .IN8(na2264_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y113     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a761_1 ( .OUT(na761_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2668_2), .IN8(na2265_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x99y114     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a762_1 ( .OUT(na762_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2266_2), .IN6(na2669_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y106     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a763_1 ( .OUT(na763_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2670_2), .IN6(na2267_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x95y87     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a764_1 ( .OUT(na764_1), .IN1(na2671_1), .IN2(na2268_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y102     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2672_2), .IN8(na2269_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y91     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a766_1 ( .OUT(na766_1), .IN1(na2673_1), .IN2(na2270_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y106     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a767_1 ( .OUT(na767_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3153_1), .IN6(na2674_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y106     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a768_1 ( .OUT(na768_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3154_2), .IN8(na2675_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y88     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a769_1 ( .OUT(na769_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2676_2), .IN8(na3155_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y112     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a770_1 ( .OUT(na770_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2677_1), .IN8(na3156_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x92y92     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a771_1 ( .OUT(na771_1), .IN1(na3157_1), .IN2(na2678_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y81     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a772_1 ( .OUT(na772_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2679_1), .IN6(na3158_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x92y95     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a773_1 ( .OUT(na773_1), .IN1(na3159_1), .IN2(na2680_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y70     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a774_1 ( .OUT(na774_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3160_2), .IN8(na2681_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y115     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2682_1), .IN6(na2271_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y103     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a776_1 ( .OUT(na776_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2272_2), .IN6(na2683_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y112     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2684_2), .IN6(na2273_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x107y114     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a778_1 ( .OUT(na778_1), .IN1(na2685_1), .IN2(na2274_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y101     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2275_1), .IN6(na2686_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x104y72     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a780_1 ( .OUT(na780_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2276_2), .IN4(na2687_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y98     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2688_2), .IN6(na2277_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y70     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a782_1 ( .OUT(na782_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2689_1), .IN6(na2278_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y109     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2690_2), .IN6(na2223_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y101     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a784_1 ( .OUT(na784_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2691_1), .IN6(na2224_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x108y109     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_1 ( .OUT(na785_1), .IN1(na2225_1), .IN2(na2692_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y111     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a786_1 ( .OUT(na786_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2226_2), .IN8(na2693_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x106y90     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1), .IN1(na2227_1), .IN2(na2694_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y68     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a788_1 ( .OUT(na788_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2228_2), .IN8(na2695_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y87     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2696_2), .IN8(na2229_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y81     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a790_1 ( .OUT(na790_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2230_2), .IN6(na2697_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y111     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_1 ( .OUT(na791_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2698_2), .IN6(na2231_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x126y106     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a792_1 ( .OUT(na792_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2232_2), .IN4(na2699_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y112     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a793_1 ( .OUT(na793_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2233_1), .IN6(na2700_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x100y113     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a794_1 ( .OUT(na794_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2234_2), .IN4(na2701_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y109     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a795_1 ( .OUT(na795_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2235_1), .IN6(na2702_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y86     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_1 ( .OUT(na796_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2703_1), .IN6(na2236_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y100     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2237_1), .IN6(na2704_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y91     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a798_1 ( .OUT(na798_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2705_1), .IN6(na2238_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y115     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a799_1 ( .OUT(na799_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3202_2), .IN7(~na800_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y115     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a800_4 ( .OUT(na800_2), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y116     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a801_1 ( .OUT(na801_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3203_1), .IN8(~na4197_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y116     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a802_4 ( .OUT(na802_2), .IN1(1'b1), .IN2(na3204_2), .IN3(~na800_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y116     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a803_1 ( .OUT(na803_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3205_1), .IN7(~na800_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y115     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a804_4 ( .OUT(na804_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na800_2), .IN4(na3206_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y113     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a805_1 ( .OUT(na805_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3207_1), .IN6(1'b1), .IN7(~na800_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y115     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a806_4 ( .OUT(na806_2), .IN1(na3208_2), .IN2(1'b1), .IN3(~na800_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y96     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a807_1 ( .OUT(na807_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na808_2), .IN6(1'b0), .IN7(na848_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x141y111     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a808_4 ( .OUT(na808_2), .IN1(1'b0), .IN2(na838_1), .IN3(na809_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y109     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na835_1), .IN6(na831_1), .IN7(na810_1), .IN8(~na834_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y111     80'h00_0018_00_0040_0A7A_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a810_1 ( .OUT(na810_1), .IN1(na811_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4206_2), .IN5(na3699_2), .IN6(~na830_1), .IN7(na815_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y115     80'h00_0018_00_0040_0AF5_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a811_1 ( .OUT(na811_1), .IN1(~na1834_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(~na3700_1), .IN6(na4399_2), .IN7(~na824_1),
                     .IN8(na1836_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x148y115     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a812_4 ( .OUT(na812_2), .IN1(na3025_1), .IN2(1'b0), .IN3(~na3019_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x147y116     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a813_1 ( .OUT(na813_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3025_2), .IN6(na3022_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y111     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a814_1 ( .OUT(na814_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3025_1), .IN6(~na4362_2), .IN7(na3021_2),
                     .IN8(na4364_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y115     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a815_4 ( .OUT(na815_2), .IN1(~na3024_1), .IN2(na3022_1), .IN3(na3023_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y116     80'h00_0060_00_0000_0C06_FF56
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a816_4 ( .OUT(na816_2), .IN1(na4202_2), .IN2(na813_1), .IN3(~na3018_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x147y111     80'h00_0018_00_0040_0C89_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1), .IN1(na3025_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na4363_2), .IN5(na3025_2), .IN6(1'b1), .IN7(na3023_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y112     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a818_1 ( .OUT(na818_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3024_1), .IN6(na3022_1), .IN7(na3019_1),
                     .IN8(na4363_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x143y114     80'h00_0018_00_0000_0666_3DED
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a819_1 ( .OUT(na819_1), .IN1(na814_1), .IN2(~na816_2), .IN3(~na815_2), .IN4(~na4199_2), .IN5(na4400_2), .IN6(~na818_1), .IN7(1'b1),
                     .IN8(na822_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x148y114     80'h00_0018_00_0000_0C66_3B00
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a822_1 ( .OUT(na822_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na823_1), .IN6(na3705_1), .IN7(1'b1), .IN8(na4361_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y113     80'h00_0018_00_0000_0C66_5A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a823_1 ( .OUT(na823_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3025_1), .IN6(1'b0), .IN7(~na3023_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y115     80'h00_0018_00_0000_0666_5A69
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a824_1 ( .OUT(na824_1), .IN1(na814_1), .IN2(~na826_2), .IN3(~na3023_2), .IN4(~na827_1), .IN5(na3707_2), .IN6(1'b0), .IN7(~na3018_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y114     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a826_4 ( .OUT(na826_2), .IN1(~na823_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3704_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y118     80'h00_0018_00_0040_0AE1_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1), .IN1(1'b1), .IN2(~na818_1), .IN3(~na815_2), .IN4(1'b1), .IN5(1'b1), .IN6(na813_1), .IN7(na3018_1),
                     .IN8(na3709_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x146y113     80'h00_0060_00_0000_0C08_FF59
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a828_4 ( .OUT(na828_2), .IN1(~na3024_1), .IN2(~na3022_1), .IN3(na812_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x147y112     80'h00_0018_00_0040_0C33_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a829_1 ( .OUT(na829_1), .IN1(~na3025_2), .IN2(~na4360_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na814_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y118     80'h00_0018_00_0040_0AF8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a830_1 ( .OUT(na830_1), .IN1(na1834_1), .IN2(1'b1), .IN3(~na824_1), .IN4(1'b1), .IN5(na4285_2), .IN6(na819_1), .IN7(na3711_1),
                     .IN8(~na1836_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y110     80'h00_0018_00_0040_0AB5_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a831_1 ( .OUT(na831_1), .IN1(1'b1), .IN2(~na833_1), .IN3(na832_1), .IN4(1'b1), .IN5(~na814_1), .IN6(na4402_2), .IN7(1'b1),
                     .IN8(na4204_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y113     80'h00_0018_00_0040_0AF5_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a832_1 ( .OUT(na832_1), .IN1(1'b1), .IN2(na819_1), .IN3(na824_1), .IN4(1'b1), .IN5(~na1834_1), .IN6(na3713_1), .IN7(~na4286_2),
                     .IN8(na1836_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y116     80'h00_0018_00_0040_0AF5_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a833_1 ( .OUT(na833_1), .IN1(1'b1), .IN2(na819_1), .IN3(1'b1), .IN4(na1836_2), .IN5(~na1834_1), .IN6(na4284_2), .IN7(~na824_1),
                     .IN8(na3714_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y108     80'h00_0018_00_0040_0A76_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a834_1 ( .OUT(na834_1), .IN1(1'b1), .IN2(na833_1), .IN3(1'b1), .IN4(na4198_2), .IN5(na814_1), .IN6(~na818_1), .IN7(~na3712_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y107     80'h00_0018_00_0040_0ADB_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a835_1 ( .OUT(na835_1), .IN1(1'b1), .IN2(~na830_1), .IN3(~na832_1), .IN4(1'b1), .IN5(~na4209_2), .IN6(1'b1), .IN7(na3716_1),
                     .IN8(~na837_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x148y107     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a836_4 ( .OUT(na836_2), .IN1(na823_1), .IN2(1'b0), .IN3(na815_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y106     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a837_1 ( .OUT(na837_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3025_2), .IN6(1'b0), .IN7(na3021_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y110     80'h00_0018_00_0000_0666_AA9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a838_1 ( .OUT(na838_1), .IN1(na840_1), .IN2(1'b0), .IN3(na3717_2), .IN4(~na841_1), .IN5(na844_1), .IN6(1'b0), .IN7(na3717_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y109     80'h00_0018_00_0040_0AD3_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a840_1 ( .OUT(na840_1), .IN1(1'b1), .IN2(na833_1), .IN3(1'b1), .IN4(~na4198_2), .IN5(~na4209_2), .IN6(1'b1), .IN7(na815_2),
                     .IN8(na4206_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y114     80'h00_0018_00_0040_0A72_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a841_1 ( .OUT(na841_1), .IN1(na811_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4208_2), .IN5(na3720_1), .IN6(~na4210_2), .IN7(na842_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x144y113     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a842_4 ( .OUT(na842_2), .IN1(na814_1), .IN2(1'b0), .IN3(~na812_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x141y113     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a843_1 ( .OUT(na843_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na813_1), .IN7(na812_2), .IN8(~na837_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y109     80'h00_0018_00_0040_0ADB_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a844_1 ( .OUT(na844_1), .IN1(1'b1), .IN2(~na830_1), .IN3(~na832_1), .IN4(1'b1), .IN5(~na847_1), .IN6(1'b1), .IN7(na3721_1),
                     .IN8(~na845_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x140y114     80'h00_0060_00_0000_0C06_FFA3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a845_4 ( .OUT(na845_2), .IN1(1'b0), .IN2(~na846_1), .IN3(na3018_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x141y116     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a846_1 ( .OUT(na846_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na823_1), .IN6(~na813_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y109     80'h00_0018_00_0000_0C66_5600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_1 ( .OUT(na847_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3025_2), .IN6(na818_1), .IN7(~na3019_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y111     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a848_1 ( .OUT(na848_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na849_1), .IN6(na850_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y113     80'h00_0018_00_0040_0AE7_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a849_1 ( .OUT(na849_1), .IN1(1'b1), .IN2(~na846_1), .IN3(1'b1), .IN4(~na4198_2), .IN5(1'b1), .IN6(~na830_1), .IN7(~na3018_1),
                     .IN8(na3722_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y110     80'h00_0018_00_0040_0AE7_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a850_1 ( .OUT(na850_1), .IN1(1'b1), .IN2(~na833_1), .IN3(~na832_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4211_2), .IN7(~na842_2),
                     .IN8(na3723_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x131y93     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a851_1 ( .OUT(na851_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3724_1), .IN4(na807_1), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y107     80'h00_0018_00_0000_0666_9639
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a852_1 ( .OUT(na852_1), .IN1(~na849_1), .IN2(na856_2), .IN3(1'b0), .IN4(~na834_1), .IN5(na835_1), .IN6(na850_1), .IN7(na853_1),
                     .IN8(~na859_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x142y109     80'h00_0018_00_0000_0666_AC9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_1 ( .OUT(na853_1), .IN1(na840_1), .IN2(1'b0), .IN3(na3717_2), .IN4(~na854_1), .IN5(1'b0), .IN6(na855_1), .IN7(na3717_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y108     80'h00_0018_00_0040_0AD8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a854_1 ( .OUT(na854_1), .IN1(na811_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4208_2), .IN5(na847_1), .IN6(1'b0), .IN7(na842_2),
                     .IN8(~na3723_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y108     80'h00_0018_00_0040_0ABC_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a855_1 ( .OUT(na855_1), .IN1(1'b1), .IN2(na830_1), .IN3(na832_1), .IN4(1'b1), .IN5(na843_1), .IN6(na3726_2), .IN7(1'b1),
                     .IN8(~na845_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y104     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a856_4 ( .OUT(na856_2), .IN1(1'b0), .IN2(na858_1), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y107     80'h00_0018_00_0040_0AD4_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_1 ( .OUT(na857_1), .IN1(na4207_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4208_2), .IN5(na847_1), .IN6(1'b0), .IN7(~na3721_1),
                     .IN8(na845_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x143y110     80'h00_0018_00_0040_0CC7_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a858_1 ( .OUT(na858_1), .IN1(na3728_2), .IN2(na846_1), .IN3(~na842_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na830_1), .IN7(1'b1),
                     .IN8(na4198_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x140y108     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a859_4 ( .OUT(na859_2), .IN1(~na844_1), .IN2(na831_1), .IN3(na810_1), .IN4(~na841_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x139y98     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a861_1 ( .OUT(na861_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na852_1), .IN6(na3729_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y94     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a862_4 ( .OUT(na862_2), .IN1(na808_2), .IN2(1'b0), .IN3(na863_2), .IN4(na864_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x138y105     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a863_4 ( .OUT(na863_2), .IN1(1'b0), .IN2(na856_2), .IN3(na853_1), .IN4(na859_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y112     80'h00_0018_00_0000_0666_9636
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a864_1 ( .OUT(na864_1), .IN1(na849_1), .IN2(na855_1), .IN3(1'b0), .IN4(~na854_1), .IN5(na835_1), .IN6(na850_1), .IN7(na809_1),
                     .IN8(~na834_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y88     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a865_1 ( .OUT(na865_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3730_1), .IN6(na862_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x136y97     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a866_4 ( .OUT(na866_2), .IN1(1'b0), .IN2(1'b0), .IN3(na867_1), .IN4(na864_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y109     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a867_1 ( .OUT(na867_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na868_2), .IN6(~na838_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y107     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a868_4 ( .OUT(na868_2), .IN1(na870_1), .IN2(~na869_1), .IN3(na4212_2), .IN4(na854_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y108     80'h00_0018_00_0040_0AE5_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1), .IN1(1'b1), .IN2(na830_1), .IN3(~na832_1), .IN4(1'b1), .IN5(1'b1), .IN6(na818_1), .IN7(~na836_2),
                     .IN8(na3731_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y105     80'h00_0018_00_0040_0AD0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_1 ( .OUT(na870_1), .IN1(na811_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4208_2), .IN5(na814_1), .IN6(1'b0), .IN7(na3732_1),
                     .IN8(na837_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y92     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_1 ( .OUT(na871_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na866_2), .IN8(na3733_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y78     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a872_1 ( .OUT(na872_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na873_1), .IN8(~na864_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x142y99     80'h00_0018_00_0000_0C66_A900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a873_1 ( .OUT(na873_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na868_2), .IN6(na856_2), .IN7(na853_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y78     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a874_1 ( .OUT(na874_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3734_2), .IN8(na872_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x127y73     80'h00_0060_00_0000_0C06_FF96
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a875_4 ( .OUT(na875_2), .IN1(na868_2), .IN2(na838_1), .IN3(na809_1), .IN4(~na4213_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y75     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a876_1 ( .OUT(na876_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na875_2), .IN6(na3735_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y91     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a877_4 ( .OUT(na877_2), .IN1(1'b0), .IN2(na879_2), .IN3(na863_2), .IN4(na878_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x132y104     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_1 ( .OUT(na878_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na868_2), .IN6(~na856_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y108     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a879_4 ( .OUT(na879_2), .IN1(na844_1), .IN2(1'b0), .IN3(1'b0), .IN4(na841_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y84     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a880_1 ( .OUT(na880_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na877_2), .IN6(na3736_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x130y83     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a881_1 ( .OUT(na881_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na870_1), .IN6(~na869_1), .IN7(na853_1), .IN8(na859_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y77     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_1 ( .OUT(na883_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na881_1), .IN8(na3737_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x142y104     80'h00_0018_00_0000_0666_09C6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a884_1 ( .OUT(na884_1), .IN1(na911_2), .IN2(na919_2), .IN3(1'b0), .IN4(na912_1), .IN5(~na913_1), .IN6(na885_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y102     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a885_4 ( .OUT(na885_2), .IN1(1'b0), .IN2(1'b0), .IN3(na886_1), .IN4(na905_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y109     80'h00_0018_00_0040_0ABD_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a886_1 ( .OUT(na886_1), .IN1(1'b1), .IN2(~na887_1), .IN3(1'b1), .IN4(na904_1), .IN5(~na903_1), .IN6(na3738_2), .IN7(1'b1),
                     .IN8(~na4365_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y100     80'h00_0018_00_0040_0AFC_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a887_1 ( .OUT(na887_1), .IN1(~na1839_1), .IN2(1'b1), .IN3(na888_1), .IN4(1'b1), .IN5(na3739_1), .IN6(na1843_2), .IN7(~na4403_2),
                     .IN8(~na1841_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x150y107     80'h00_0018_00_0000_0666_96C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a888_1 ( .OUT(na888_1), .IN1(~na3027_1), .IN2(1'b0), .IN3(1'b0), .IN4(na893_2), .IN5(na3741_2), .IN6(na4370_2), .IN7(~na889_1),
                     .IN8(na896_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x146y107     80'h00_0018_00_0000_0C66_EC00
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a889_1 ( .OUT(na889_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na890_2), .IN7(~na3742_1), .IN8(~na893_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x149y106     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a890_4 ( .OUT(na890_2), .IN1(na892_2), .IN2(na3744_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y110     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3030_1), .IN8(~na3033_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x147y103     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a892_4 ( .OUT(na892_2), .IN1(~na4369_2), .IN2(na3029_2), .IN3(na4372_2), .IN4(~na3031_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y110     80'h00_0060_00_0000_0C06_FF9A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a893_4 ( .OUT(na893_2), .IN1(na4367_2), .IN2(1'b0), .IN3(na3030_1), .IN4(~na3032_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x147y110     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a894_4 ( .OUT(na894_2), .IN1(na4220_2), .IN2(1'b0), .IN3(na3026_2), .IN4(na891_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x148y98     80'h00_0018_00_0040_0C89_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a896_1 ( .OUT(na896_1), .IN1(na4369_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na3033_1), .IN5(na4367_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na3033_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y103     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3027_1), .IN6(na4370_2), .IN7(na3030_1), .IN8(~na3032_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x147y105     80'h00_0018_00_0000_0C88_56FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a899_1 ( .OUT(na899_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3027_1), .IN6(~na4371_2), .IN7(na900_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y105     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_1 ( .OUT(na900_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4369_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na3031_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x146y101     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a901_1 ( .OUT(na901_1), .IN1(na892_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3027_1), .IN6(~na4371_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x141y106     80'h00_0018_00_0000_0C88_96FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a902_1 ( .OUT(na902_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3027_1), .IN6(na4370_2), .IN7(na3030_1),
                     .IN8(na3032_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y103     80'h00_0018_00_0040_0AF3_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a903_1 ( .OUT(na903_1), .IN1(1'b1), .IN2(~na4289_2), .IN3(~na888_1), .IN4(1'b1), .IN5(~na1839_1), .IN6(~na1843_2), .IN7(na4290_2),
                     .IN8(na3749_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y100     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a904_1 ( .OUT(na904_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na900_1), .IN8(~na891_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x146y98     80'h00_0018_00_0040_0C7E_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a905_1 ( .OUT(na905_1), .IN1(1'b1), .IN2(~na4225_2), .IN3(~na909_2), .IN4(na3750_2), .IN5(~na4224_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y104     80'h00_0018_00_0040_0AF6_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a906_1 ( .OUT(na906_1), .IN1(1'b1), .IN2(na1843_2), .IN3(1'b1), .IN4(~na1841_1), .IN5(na1839_1), .IN6(~na4287_2), .IN7(~na888_1),
                     .IN8(na3751_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y100     80'h00_0018_00_0040_0AF1_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a907_1 ( .OUT(na907_1), .IN1(1'b1), .IN2(na1843_2), .IN3(1'b1), .IN4(na4288_2), .IN5(~na4217_2), .IN6(na3752_2), .IN7(na888_1),
                     .IN8(na1841_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x147y99     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a908_1 ( .OUT(na908_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na892_2), .IN6(1'b0), .IN7(na4366_2), .IN8(na3033_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y99     80'h00_0060_00_0000_0C06_FF65
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a909_4 ( .OUT(na909_2), .IN1(~na3027_1), .IN2(1'b0), .IN3(na897_1), .IN4(na3033_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x141y101     80'h00_0060_00_0000_0C06_FFE7
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a911_4 ( .OUT(na911_2), .IN1(na892_2), .IN2(na4222_2), .IN3(~na897_1), .IN4(~na906_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x144y100     80'h00_0018_00_0040_0CA7_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a912_1 ( .OUT(na912_1), .IN1(na4219_2), .IN2(~na924_1), .IN3(na900_1), .IN4(1'b1), .IN5(1'b1), .IN6(na887_1), .IN7(1'b1),
                     .IN8(~na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y105     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a913_1 ( .OUT(na913_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na917_1), .IN6(1'b0), .IN7(1'b0), .IN8(na914_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y98     80'h00_0018_00_0040_0AD0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a914_1 ( .OUT(na914_1), .IN1(1'b1), .IN2(na887_1), .IN3(~na915_1), .IN4(1'b1), .IN5(na908_1), .IN6(1'b0), .IN7(na3756_1),
                     .IN8(na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y101     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a915_1 ( .OUT(na915_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3027_1), .IN6(~na4370_2), .IN7(na4218_2),
                     .IN8(na916_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y104     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a916_1 ( .OUT(na916_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3029_2), .IN7(1'b0), .IN8(na3033_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y97     80'h00_0018_00_0040_0A7E_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a917_1 ( .OUT(na917_1), .IN1(~na903_1), .IN2(1'b1), .IN3(1'b1), .IN4(na906_1), .IN5(na3757_2), .IN6(~na918_2), .IN7(~na909_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y98     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a918_4 ( .OUT(na918_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3026_2), .IN4(~na904_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x141y100     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a919_4 ( .OUT(na919_2), .IN1(na920_1), .IN2(na921_1), .IN3(~na922_1), .IN4(~na923_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y103     80'h00_0018_00_0040_0AB5_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_1 ( .OUT(na920_1), .IN1(1'b1), .IN2(~na887_1), .IN3(na900_1), .IN4(1'b1), .IN5(~na903_1), .IN6(na3758_1), .IN7(1'b1),
                     .IN8(na893_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y98     80'h00_0018_00_0040_0ADB_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a921_1 ( .OUT(na921_1), .IN1(na4224_2), .IN2(1'b1), .IN3(~na897_1), .IN4(1'b1), .IN5(~na892_2), .IN6(1'b1), .IN7(na3759_2),
                     .IN8(~na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y101     80'h00_0018_00_0040_0ABC_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a922_1 ( .OUT(na922_1), .IN1(na892_2), .IN2(1'b1), .IN3(na897_1), .IN4(1'b1), .IN5(na3760_1), .IN6(na887_1), .IN7(1'b1),
                     .IN8(~na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y102     80'h00_0018_00_0040_0ADB_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a923_1 ( .OUT(na923_1), .IN1(~na903_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na906_1), .IN5(~na4228_2), .IN6(1'b1), .IN7(na3761_2),
                     .IN8(~na916_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y104     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a924_1 ( .OUT(na924_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na900_1), .IN8(na893_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x136y96     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a925_1 ( .OUT(na925_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3762_2), .IN8(na884_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y100     80'h00_0018_00_0000_0666_9A66
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a926_1 ( .OUT(na926_1), .IN1(na931_1), .IN2(na885_2), .IN3(~na928_1), .IN4(~na923_1), .IN5(na911_2), .IN6(1'b0), .IN7(~na922_1),
                     .IN8(na912_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y95     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a928_1 ( .OUT(na928_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na920_1), .IN6(na921_1), .IN7(~na929_1), .IN8(na930_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x142y95     80'h00_0018_00_0040_0C17_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a929_1 ( .OUT(na929_1), .IN1(~na3757_2), .IN2(na918_2), .IN3(na909_2), .IN4(1'b0), .IN5(na4224_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x142y96     80'h00_0018_00_0040_0C5B_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a930_1 ( .OUT(na930_1), .IN1(~na908_1), .IN2(na3764_1), .IN3(1'b1), .IN4(na904_1), .IN5(1'b1), .IN6(~na887_1), .IN7(1'b1),
                     .IN8(~na4223_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y97     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a931_1 ( .OUT(na931_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na917_1), .IN6(~na933_1), .IN7(~na932_1), .IN8(na914_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x142y97     80'h00_0018_00_0040_0CCB_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a932_1 ( .OUT(na932_1), .IN1(na3760_1), .IN2(na887_1), .IN3(1'b1), .IN4(~na907_1), .IN5(na908_1), .IN6(1'b1), .IN7(~na909_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y98     80'h00_0018_00_0040_0AE3_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a933_1 ( .OUT(na933_1), .IN1(na903_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na906_1), .IN5(1'b1), .IN6(~na918_2), .IN7(na915_1),
                     .IN8(na3766_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x133y93     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a934_1 ( .OUT(na934_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3767_2), .IN4(na926_1), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y84     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a935_1 ( .OUT(na935_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na937_2), .IN7(~na938_1), .IN8(na936_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y104     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a936_1 ( .OUT(na936_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na913_1), .IN6(na919_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y92     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a937_4 ( .OUT(na937_2), .IN1(na931_1), .IN2(1'b0), .IN3(na928_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y99     80'h00_0018_00_0000_0666_3999
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a938_1 ( .OUT(na938_1), .IN1(~na939_2), .IN2(na885_2), .IN3(~na922_1), .IN4(na912_1), .IN5(~na911_2), .IN6(na919_2), .IN7(1'b0),
                     .IN8(~na923_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x141y97     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a939_4 ( .OUT(na939_2), .IN1(na911_2), .IN2(~na933_1), .IN3(~na932_1), .IN4(na912_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x133y81     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a940_1 ( .OUT(na940_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3768_1), .IN4(na935_1), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y95     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a941_1 ( .OUT(na941_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na943_2), .IN7(na938_1), .IN8(na942_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x138y104     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a942_4 ( .OUT(na942_2), .IN1(na913_1), .IN2(~na919_2), .IN3(na4226_2), .IN4(na912_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y102     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a943_4 ( .OUT(na943_2), .IN1(na4227_2), .IN2(na944_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y96     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a944_4 ( .OUT(na944_2), .IN1(na4230_2), .IN2(~na945_1), .IN3(na932_1), .IN4(~na946_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y102     80'h00_0018_00_0040_0A74_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_1 ( .OUT(na945_1), .IN1(~na903_1), .IN2(1'b1), .IN3(1'b1), .IN4(na906_1), .IN5(na3769_2), .IN6(na924_1), .IN7(~na897_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x142y98     80'h00_0018_00_0040_0CBD_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a946_1 ( .OUT(na946_1), .IN1(~na892_2), .IN2(1'b1), .IN3(na3770_2), .IN4(~na916_1), .IN5(1'b1), .IN6(na887_1), .IN7(1'b1),
                     .IN8(na907_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y92     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a947_1 ( .OUT(na947_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na941_1), .IN8(na3771_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x134y70     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a948_4 ( .OUT(na948_2), .IN1(1'b0), .IN2(1'b0), .IN3(na938_1), .IN4(na949_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y82     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a949_4 ( .OUT(na949_2), .IN1(na939_2), .IN2(~na944_2), .IN3(na929_1), .IN4(na930_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y72     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a951_1 ( .OUT(na951_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3772_1), .IN8(na948_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x128y65     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a952_4 ( .OUT(na952_2), .IN1(1'b0), .IN2(1'b0), .IN3(na953_1), .IN4(~na949_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x128y73     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a953_1 ( .OUT(na953_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na931_1), .IN6(~na919_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y67     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a954_1 ( .OUT(na954_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na952_2), .IN8(na3773_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y80     80'h00_0018_00_0000_0666_A066
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a955_1 ( .OUT(na955_1), .IN1(~na939_2), .IN2(~na944_2), .IN3(na929_1), .IN4(na930_1), .IN5(1'b0), .IN6(1'b0), .IN7(na928_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y76     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a956_1 ( .OUT(na956_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3774_2), .IN8(na955_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y67     80'h00_0060_00_0000_0C06_FFC3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a957_4 ( .OUT(na957_2), .IN1(1'b0), .IN2(~na937_2), .IN3(1'b0), .IN4(na949_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y71     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a958_1 ( .OUT(na958_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na957_2), .IN6(na3775_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y105     80'h00_0018_00_0000_0666_A636
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a959_1 ( .OUT(na959_1), .IN1(~na987_1), .IN2(~na985_1), .IN3(1'b0), .IN4(~na996_2), .IN5(na990_1), .IN6(na961_1), .IN7(na982_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x135y112     80'h00_0018_00_0000_0C66_E7FF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a961_1 ( .OUT(na961_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na963_2), .IN6(na962_1), .IN7(~na981_1), .IN8(~na969_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y118     80'h00_0018_00_0040_0AF8_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a962_1 ( .OUT(na962_1), .IN1(1'b1), .IN2(na4291_2), .IN3(~na4241_2), .IN4(1'b1), .IN5(na4293_2), .IN6(na970_1), .IN7(na3778_2),
                     .IN8(~na1848_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y115     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a963_4 ( .OUT(na963_2), .IN1(~na3039_2), .IN2(na4378_2), .IN3(na3037_2), .IN4(~na3041_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y116     80'h00_0018_00_0000_0C66_3C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a964_1 ( .OUT(na964_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3038_1), .IN7(1'b0), .IN8(~na3041_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x138y115     80'h00_0060_00_0000_0C06_FFC3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a965_4 ( .OUT(na965_2), .IN1(1'b0), .IN2(~na3035_1), .IN3(1'b0), .IN4(na3041_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x138y113     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a966_4 ( .OUT(na966_2), .IN1(~na3040_1), .IN2(na3038_1), .IN3(na4376_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x137y116     80'h00_0018_00_0000_0C66_A900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a967_1 ( .OUT(na967_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3034_2), .IN6(na964_1), .IN7(na966_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x142y116     80'h00_0018_00_0040_0C89_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a968_1 ( .OUT(na968_1), .IN1(na4377_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na3041_1), .IN5(na3039_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na3041_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y114     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a969_1 ( .OUT(na969_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3040_1), .IN6(na3035_1), .IN7(na4374_2),
                     .IN8(na3041_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x135y116     80'h00_0018_00_0000_0666_D3ED
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a970_1 ( .OUT(na970_1), .IN1(na963_2), .IN2(~na967_1), .IN3(~na966_2), .IN4(~na4235_2), .IN5(1'b1), .IN6(na973_1), .IN7(na4404_2),
                     .IN8(~na969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x141y114     80'h00_0018_00_0000_0C66_3D00
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_1 ( .OUT(na973_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3782_2), .IN6(~na974_1), .IN7(1'b1), .IN8(na4375_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y114     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a974_1 ( .OUT(na974_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3039_2), .IN6(1'b0), .IN7(1'b0), .IN8(na3041_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y115     80'h00_0018_00_0000_0666_65A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a975_1 ( .OUT(na975_1), .IN1(~na3034_2), .IN2(~na977_1), .IN3(na3784_1), .IN4(1'b0), .IN5(~na3039_2), .IN6(1'b0), .IN7(na978_2),
                     .IN8(na4232_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y114     80'h00_0018_00_0040_0AB9_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a977_1 ( .OUT(na977_1), .IN1(1'b1), .IN2(~na964_1), .IN3(na966_2), .IN4(1'b1), .IN5(~na3034_2), .IN6(na3785_2), .IN7(1'b0),
                     .IN8(~na969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y115     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a978_4 ( .OUT(na978_2), .IN1(1'b1), .IN2(~na974_1), .IN3(1'b1), .IN4(na3781_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x136y112     80'h00_0018_00_0000_0C88_59FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a979_1 ( .OUT(na979_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3040_1), .IN6(~na3038_1), .IN7(na965_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x137y113     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a980_1 ( .OUT(na980_1), .IN1(na963_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4373_2), .IN8(~na3041_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y117     80'h00_0018_00_0040_0AFC_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a981_1 ( .OUT(na981_1), .IN1(na975_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4238_2), .IN5(na3788_2), .IN6(na4294_2), .IN7(~na1846_2),
                     .IN8(~na1848_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x126y113     80'h00_0018_00_0040_0C3D_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a982_1 ( .OUT(na982_1), .IN1(~na1001_2), .IN2(1'b1), .IN3(na966_2), .IN4(na4239_2), .IN5(1'b1), .IN6(~na984_1), .IN7(1'b1),
                     .IN8(~na983_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y116     80'h00_0018_00_0040_0AF3_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a983_1 ( .OUT(na983_1), .IN1(1'b1), .IN2(na970_1), .IN3(~na1846_2), .IN4(1'b1), .IN5(~na4405_2), .IN6(~na4240_2), .IN7(na3790_1),
                     .IN8(na1848_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y116     80'h00_0018_00_0040_0AF8_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a984_1 ( .OUT(na984_1), .IN1(1'b1), .IN2(na970_1), .IN3(1'b1), .IN4(~na1848_1), .IN5(na975_1), .IN6(na3792_2), .IN7(na1846_2),
                     .IN8(~na4292_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y112     80'h00_0018_00_0040_0AB7_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a985_1 ( .OUT(na985_1), .IN1(1'b1), .IN2(na962_1), .IN3(1'b1), .IN4(na983_1), .IN5(~na3034_2), .IN6(~na995_2), .IN7(1'b1),
                     .IN8(na986_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y116     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a986_4 ( .OUT(na986_2), .IN1(na4233_2), .IN2(~na974_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x127y113     80'h00_0018_00_0040_0CE7_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a987_1 ( .OUT(na987_1), .IN1(na3794_1), .IN2(~na4244_2), .IN3(~na989_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na984_1), .IN7(na981_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y115     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a988_1 ( .OUT(na988_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na963_2), .IN6(1'b0), .IN7(na965_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x132y113     80'h00_0060_00_0000_0C06_FFC9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a989_4 ( .OUT(na989_2), .IN1(na4237_2), .IN2(~na3035_1), .IN3(1'b0), .IN4(na3041_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y109     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a990_1 ( .OUT(na990_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na991_1), .IN7(1'b0), .IN8(na994_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y118     80'h00_0018_00_0040_0A70_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a991_1 ( .OUT(na991_1), .IN1(na4242_2), .IN2(1'b1), .IN3(na992_2), .IN4(1'b1), .IN5(na3795_1), .IN6(na984_1), .IN7(na4245_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x134y117     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a992_4 ( .OUT(na992_2), .IN1(1'b0), .IN2(na964_1), .IN3(~na965_2), .IN4(na993_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y114     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a993_1 ( .OUT(na993_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3037_2), .IN8(na3041_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y116     80'h00_0018_00_0040_0A7E_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a994_1 ( .OUT(na994_1), .IN1(1'b1), .IN2(~na962_1), .IN3(na981_1), .IN4(1'b1), .IN5(na4406_2), .IN6(~na995_2), .IN7(~na989_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y116     80'h00_0060_00_0000_0C06_FF3A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a995_4 ( .OUT(na995_2), .IN1(na3034_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na986_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x132y112     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a996_4 ( .OUT(na996_2), .IN1(na998_1), .IN2(~na999_1), .IN3(~na1000_1), .IN4(na997_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y110     80'h00_0018_00_0040_0AE9_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a997_1 ( .OUT(na997_1), .IN1(1'b1), .IN2(na962_1), .IN3(1'b1), .IN4(~na983_1), .IN5(1'b1), .IN6(na974_1), .IN7(na966_2),
                     .IN8(~na4250_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y111     80'h00_0018_00_0040_0ABD_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a998_1 ( .OUT(na998_1), .IN1(~na4237_2), .IN2(1'b1), .IN3(na981_1), .IN4(1'b1), .IN5(~na963_2), .IN6(na3798_1), .IN7(1'b1),
                     .IN8(~na4243_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y114     80'h00_0018_00_0040_0AE3_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_1 ( .OUT(na999_1), .IN1(na963_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na969_1), .IN5(1'b1), .IN6(~na984_1), .IN7(na3799_2),
                     .IN8(na983_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y113     80'h00_0018_00_0040_0ADB_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1), .IN1(1'b1), .IN2(~na962_1), .IN3(~na981_1), .IN4(1'b1), .IN5(~na1001_2), .IN6(1'b1), .IN7(na3800_1),
                      .IN8(~na993_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x133y113     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1001_4 ( .OUT(na1001_2), .IN1(1'b0), .IN2(na974_1), .IN3(na966_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y96     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1002_1 ( .OUT(na1002_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na959_1), .IN6(na3801_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y110     80'h00_0018_00_0000_0666_5699
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_1 ( .OUT(na1003_1), .IN1(na990_1), .IN2(~na999_1), .IN3(~na1005_1), .IN4(na1008_2), .IN5(na987_1), .IN6(na985_1), .IN7(~na1000_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x132y111     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1005_1 ( .OUT(na1005_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1006_1), .IN6(na961_1), .IN7(na982_1), .IN8(~na1007_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x127y115     80'h00_0018_00_0040_0C3E_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1006_1 ( .OUT(na1006_1), .IN1(1'b1), .IN2(~na984_1), .IN3(na3799_2), .IN4(na983_1), .IN5(na988_1), .IN6(1'b1), .IN7(na989_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y116     80'h00_0018_00_0040_0AE3_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1007_1 ( .OUT(na1007_1), .IN1(1'b1), .IN2(na962_1), .IN3(~na981_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na995_2), .IN7(na992_2),
                      .IN8(na3803_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x134y110     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1008_4 ( .OUT(na1008_2), .IN1(~na1009_1), .IN2(na4249_2), .IN3(na1010_1), .IN4(na997_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x133y111     80'h00_0018_00_0040_0C8E_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1), .IN1(1'b0), .IN2(na995_2), .IN3(na989_2), .IN4(~na3796_2), .IN5(1'b1), .IN6(na984_1), .IN7(~na981_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y111     80'h00_0018_00_0040_0AD3_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_1 ( .OUT(na1010_1), .IN1(1'b1), .IN2(~na962_1), .IN3(1'b1), .IN4(~na983_1), .IN5(~na988_1), .IN6(1'b1), .IN7(na3805_2),
                      .IN8(na986_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y97     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1011_1 ( .OUT(na1011_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3806_1), .IN8(na1003_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y97     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_1 ( .OUT(na1012_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1014_2), .IN7(~na1016_1), .IN8(na1013_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y110     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1013_4 ( .OUT(na1013_2), .IN1(na990_1), .IN2(1'b0), .IN3(na1005_1), .IN4(na1008_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x113y110     80'h00_0060_00_0000_0C06_FF9A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1014_4 ( .OUT(na1014_2), .IN1(na990_1), .IN2(1'b0), .IN3(~na4247_2), .IN4(na1015_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y114     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1015_1 ( .OUT(na1015_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na961_1), .IN7(na982_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y111     80'h00_0018_00_0000_0666_69A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_1 ( .OUT(na1016_1), .IN1(~na987_1), .IN2(na961_1), .IN3(na1005_1), .IN4(1'b0), .IN5(na998_1), .IN6(~na985_1), .IN7(na982_1),
                      .IN8(na997_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y90     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_1 ( .OUT(na1018_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1012_1), .IN6(na3807_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y100     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1019_4 ( .OUT(na1019_2), .IN1(1'b0), .IN2(na1020_1), .IN3(na1016_1), .IN4(~na996_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y116     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1020_1 ( .OUT(na1020_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na990_1), .IN6(~na1021_1), .IN7(~na4248_2),
                      .IN8(na1015_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y110     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1021_1 ( .OUT(na1021_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1006_1), .IN6(~na1022_1), .IN7(~na1023_1),
                      .IN8(na1007_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x129y114     80'h00_0018_00_0040_0AB8_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_1 ( .OUT(na1022_1), .IN1(1'b1), .IN2(na962_1), .IN3(na981_1), .IN4(1'b1), .IN5(na1001_2), .IN6(na3808_1), .IN7(1'b0),
                      .IN8(~na969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y115     80'h00_0018_00_0040_0CDB_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_1 ( .OUT(na1023_1), .IN1(~na963_2), .IN2(na3809_2), .IN3(1'b1), .IN4(~na993_1), .IN5(1'b1), .IN6(na984_1), .IN7(1'b1),
                      .IN8(na983_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y98     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1024_1 ( .OUT(na1024_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3810_1), .IN8(na1019_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y87     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1026_2), .IN6(1'b0), .IN7(na1016_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x117y111     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1026_4 ( .OUT(na1026_2), .IN1(na1009_1), .IN2(~na1021_1), .IN3(na1010_1), .IN4(na4252_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y83     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1025_1), .IN6(na3811_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y82     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1029_1 ( .OUT(na1029_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1014_2), .IN7(na1030_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x106y105     80'h00_0018_00_0000_0C66_A900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1009_1), .IN6(na1021_1), .IN7(na1010_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y77     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1031_1 ( .OUT(na1031_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3812_1), .IN8(na1029_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x116y106     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1032_1 ( .OUT(na1032_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na998_1), .IN6(~na1021_1), .IN7(na1005_1),
                      .IN8(na997_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y91     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3813_2), .IN8(na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x124y92     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1034_4 ( .OUT(na1034_2), .IN1(1'b0), .IN2(na1035_1), .IN3(na1030_1), .IN4(na1015_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x109y108     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_1 ( .OUT(na1035_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na990_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1008_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x113y82     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1036_1 ( .OUT(na1036_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3814_1), .IN4(na1034_2), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y87     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1037_1 ( .OUT(na1037_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3724_1), .IN8(na807_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x140y98     80'h00_0018_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1038_1 ( .OUT(na1038_1), .IN1(na852_1), .IN2(na3729_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x139y90     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3730_1), .IN6(na862_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x129y87     80'h00_0018_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1040_1 ( .OUT(na1040_1), .IN1(1'b0), .IN2(1'b0), .IN3(na866_2), .IN4(na3733_1), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x139y74     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1041_1 ( .OUT(na1041_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3734_2), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y71     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1042_1 ( .OUT(na1042_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na875_2), .IN6(na3735_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x141y83     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1043_1 ( .OUT(na1043_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na877_2), .IN6(na3736_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y76     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1044_1 ( .OUT(na1044_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na881_1), .IN8(na3737_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x140y94     80'h00_0018_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1045_1 ( .OUT(na1045_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3762_2), .IN4(na884_1), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x139y92     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1046_1 ( .OUT(na1046_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3767_2), .IN8(na926_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x139y78     80'h00_0018_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1047_1 ( .OUT(na1047_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3768_1), .IN4(na935_1), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x139y87     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1048_1 ( .OUT(na1048_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na941_1), .IN8(na3771_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y71     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1049_1 ( .OUT(na1049_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3772_1), .IN8(na948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y68     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1050_1 ( .OUT(na1050_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na952_2), .IN8(na3773_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y69     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_1 ( .OUT(na1051_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3774_2), .IN8(na955_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x135y70     80'h00_0018_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1052_1 ( .OUT(na1052_1), .IN1(na957_2), .IN2(na3775_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y98     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1053_1 ( .OUT(na1053_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na959_1), .IN6(na3801_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x131y99     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1054_1 ( .OUT(na1054_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3806_1), .IN4(na1003_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y90     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_1 ( .OUT(na1055_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1012_1), .IN6(na3807_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y93     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1056_1 ( .OUT(na1056_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3810_1), .IN8(na1019_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y83     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1057_1 ( .OUT(na1057_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1025_1), .IN6(na3811_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y78     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1058_1 ( .OUT(na1058_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3812_1), .IN8(na1029_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x120y92     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_1 ( .OUT(na1059_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3813_2), .IN4(na1032_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y84     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1060_1 ( .OUT(na1060_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3814_1), .IN8(na1034_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x133y94     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_1 ( .OUT(na1061_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3724_1), .IN4(na807_1), .IN5(1'b1), .IN6(~na16_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x138y95     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1062_1 ( .OUT(na1062_1), .IN1(1'b1), .IN2(na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(na852_1), .IN6(na3729_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x137y85     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_1 ( .OUT(na1063_1), .IN1(1'b1), .IN2(~na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3730_1), .IN6(na862_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y87     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1), .IN1(1'b1), .IN2(na16_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na866_2), .IN8(na3733_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y76     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1065_1 ( .OUT(na1065_1), .IN1(1'b1), .IN2(~na16_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3734_2), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x125y76     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1066_1 ( .OUT(na1066_1), .IN1(na875_2), .IN2(na3735_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na16_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x133y84     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1067_1 ( .OUT(na1067_1), .IN1(1'b1), .IN2(na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(na877_2), .IN6(na3736_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x129y79     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1068_1 ( .OUT(na1068_1), .IN1(1'b0), .IN2(1'b0), .IN3(na881_1), .IN4(na3737_1), .IN5(1'b1), .IN6(na16_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x133y96     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_1 ( .OUT(na1069_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3762_2), .IN8(na884_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y94     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3767_2), .IN8(na926_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y83     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_1 ( .OUT(na1071_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3768_1), .IN8(na935_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y91     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1072_1 ( .OUT(na1072_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na941_1), .IN8(na3771_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x130y74     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1073_1 ( .OUT(na1073_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3772_1), .IN4(na948_2), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y71     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1074_1 ( .OUT(na1074_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na952_2), .IN8(na3773_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x129y78     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1075_1 ( .OUT(na1075_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3774_2), .IN4(na955_1), .IN5(1'b1), .IN6(~na543_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y76     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1076_1 ( .OUT(na1076_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na957_2), .IN6(na3775_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y95     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1077_1 ( .OUT(na1077_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na959_1), .IN6(na3801_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y92     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1078_1 ( .OUT(na1078_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3806_1), .IN8(na1003_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y94     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_1 ( .OUT(na1079_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1012_1), .IN6(na3807_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x127y91     80'h00_0018_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1080_1 ( .OUT(na1080_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3810_1), .IN4(na1019_2), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x133y82     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1025_1), .IN6(na3811_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x125y78     80'h00_0018_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1082_1 ( .OUT(na1082_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3812_1), .IN4(na1029_1), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y89     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_1 ( .OUT(na1083_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3813_2), .IN8(na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y85     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1084_1 ( .OUT(na1084_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3814_1), .IN8(na1034_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y91     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_1 ( .OUT(na1085_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na19_1), .IN5(na4407_2), .IN6(1'b0), .IN7(na215_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y95     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1086_1 ( .OUT(na1086_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(1'b0), .IN6(na4408_2), .IN7(1'b0), .IN8(na263_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x119y82     80'h00_0018_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_1 ( .OUT(na1087_1), .IN1(1'b0), .IN2(na4409_2), .IN3(1'b0), .IN4(na275_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na19_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y96     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1088_1 ( .OUT(na1088_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na19_1), .IN5(na3866_1), .IN6(1'b0), .IN7(na281_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x116y80     80'h00_0018_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1089_1 ( .OUT(na1089_1), .IN1(na3867_2), .IN2(1'b0), .IN3(na293_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na19_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y85     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1090_1 ( .OUT(na1090_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na19_1), .IN5(na4412_2), .IN6(1'b0), .IN7(na298_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y89     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1091_1 ( .OUT(na1091_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na19_1), .IN5(na308_1), .IN6(1'b0), .IN7(na3869_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y82     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1092_1 ( .OUT(na1092_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na19_1), .IN5(na312_1), .IN6(1'b0), .IN7(na4414_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y94     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1093_1 ( .OUT(na1093_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3724_1), .IN8(na807_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x135y96     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1094_1 ( .OUT(na1094_1), .IN1(na852_1), .IN2(na3729_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na543_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y87     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1095_1 ( .OUT(na1095_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3730_1), .IN6(na862_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x125y92     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1096_1 ( .OUT(na1096_1), .IN1(1'b0), .IN2(1'b0), .IN3(na866_2), .IN4(na3733_1), .IN5(1'b1), .IN6(na543_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y80     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1097_1 ( .OUT(na1097_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3734_2), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y75     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1098_1 ( .OUT(na1098_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na875_2), .IN6(na3735_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y86     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1099_1 ( .OUT(na1099_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na877_2), .IN6(na3736_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y80     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1100_1 ( .OUT(na1100_1), .IN1(1'b1), .IN2(na543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na881_1), .IN8(na3737_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x138y93     80'h00_0018_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1101_1 ( .OUT(na1101_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3762_2), .IN4(na884_1), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x137y94     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1102_1 ( .OUT(na1102_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3767_2), .IN8(na926_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x137y80     80'h00_0018_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1103_1 ( .OUT(na1103_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3768_1), .IN4(na935_1), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x139y88     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1104_1 ( .OUT(na1104_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na941_1), .IN8(na3771_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y71     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1105_1 ( .OUT(na1105_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3772_1), .IN8(na948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y68     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1106_1 ( .OUT(na1106_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na952_2), .IN8(na3773_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x133y73     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1107_1 ( .OUT(na1107_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3774_2), .IN8(na955_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x132y72     80'h00_0018_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1108_1 ( .OUT(na1108_1), .IN1(na957_2), .IN2(na3775_1), .IN3(1'b0), .IN4(1'b0), .IN5(na21_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y95     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1109_1 ( .OUT(na1109_1), .IN1(1'b1), .IN2(~na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(na959_1), .IN6(na3801_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x134y96     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1110_1 ( .OUT(na1110_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3806_1), .IN4(na1003_1), .IN5(1'b1), .IN6(na16_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y87     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_1 ( .OUT(na1111_1), .IN1(1'b1), .IN2(~na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1012_1), .IN6(na3807_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y90     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1112_1 ( .OUT(na1112_1), .IN1(1'b1), .IN2(na16_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3810_1), .IN8(na1019_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y80     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1113_1 ( .OUT(na1113_1), .IN1(1'b1), .IN2(~na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1025_1), .IN6(na3811_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y77     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1114_1 ( .OUT(na1114_1), .IN1(1'b1), .IN2(na16_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3812_1), .IN8(na1029_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x122y88     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1115_1 ( .OUT(na1115_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3813_2), .IN4(na1032_1), .IN5(1'b1), .IN6(na16_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y81     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_1 ( .OUT(na1116_1), .IN1(1'b1), .IN2(na16_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3814_1), .IN8(na1034_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x120y87     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1117_1 ( .OUT(na1117_1), .IN1(1'b0), .IN2(1'b0), .IN3(na215_2), .IN4(na3863_2), .IN5(1'b1), .IN6(na57_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y89     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1118_1 ( .OUT(na1118_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3864_1), .IN8(na263_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y81     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1119_1 ( .OUT(na1119_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3865_2), .IN8(na275_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y88     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1120_1 ( .OUT(na1120_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na281_1), .IN8(na4410_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y76     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_1 ( .OUT(na1121_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na293_1), .IN8(na4411_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x115y75     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1122_1 ( .OUT(na1122_1), .IN1(1'b0), .IN2(1'b0), .IN3(na298_1), .IN4(na3868_1), .IN5(1'b1), .IN6(na57_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y82     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1123_1 ( .OUT(na1123_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(na4413_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x115y76     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1124_1 ( .OUT(na1124_1), .IN1(na312_1), .IN2(na3870_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na57_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y82     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1125_1 ( .OUT(na1125_1), .IN1(1'b1), .IN2(na1126_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na215_2), .IN8(na3863_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y72     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1126_4 ( .OUT(na1126_2), .IN1(na2415_2), .IN2(na2416_1), .IN3(na2417_1), .IN4(~na4310_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y88     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1127_1 ( .OUT(na1127_1), .IN1(1'b1), .IN2(~na1126_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3864_1), .IN8(na263_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y73     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1128_1 ( .OUT(na1128_1), .IN1(1'b1), .IN2(~na1126_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3865_2), .IN8(na275_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y88     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1), .IN1(1'b1), .IN2(na1126_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na281_1), .IN8(na4410_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y72     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1130_1 ( .OUT(na1130_1), .IN1(1'b1), .IN2(na1126_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na293_1), .IN8(na4411_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y73     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1), .IN1(1'b1), .IN2(na1126_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na298_1), .IN8(na3868_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y78     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1132_1 ( .OUT(na1132_1), .IN1(1'b1), .IN2(na1126_2), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(na4413_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1133_1 ( .OUT(na1133_1), .IN1(1'b1), .IN2(na1126_2), .IN3(1'b0), .IN4(1'b0), .IN5(na312_1), .IN6(na3870_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y89     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na539_2), .IN7(1'b1), .IN8(na1946_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x125y100     80'h00_0018_00_0040_0C4C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1137_1), .IN4(na3863_2), .IN5(1'b1), .IN6(~na1136_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x135y98     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1136_4 ( .OUT(na1136_2), .IN1(1'b0), .IN2(na3285_2), .IN3(na3151_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y101     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2450_2), .IN6(~na4311_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x121y101     80'h00_0018_00_0040_0C8C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1138_1 ( .OUT(na1138_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3864_1), .IN4(~na1139_1), .IN5(1'b1), .IN6(na1136_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y102     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2451_1), .IN8(~na4313_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y94     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3865_2), .IN8(~na1141_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y94     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4310_2), .IN5(~na2420_2), .IN6(1'b0), .IN7(~na2452_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y100     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1142_1 ( .OUT(na1142_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3866_1), .IN6(~na1143_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x109y100     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1143_1 ( .OUT(na1143_1), .IN1(~na2421_1), .IN2(~na4322_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2416_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y93     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1144_1 ( .OUT(na1144_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3867_2), .IN6(~na1145_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x115y92     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_1 ( .OUT(na1145_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4315_2), .IN4(~na2454_1), .IN5(1'b1), .IN6(na2416_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y94     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1146_1 ( .OUT(na1146_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1147_1), .IN8(na3868_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y89     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2455_2), .IN8(~na4316_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y102     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1148_1 ( .OUT(na1148_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3869_1), .IN8(~na1149_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y94     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1149_1 ( .OUT(na1149_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(~na2456_1), .IN7(1'b0), .IN8(~na2424_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x122y93     80'h00_0018_00_0040_0C13_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1150_1 ( .OUT(na1150_1), .IN1(~na1151_1), .IN2(na3870_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1136_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y85     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_1 ( .OUT(na1151_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2425_2), .IN6(~na2457_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x142y103     80'h00_0018_00_0040_0C8C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1152_1 ( .OUT(na1152_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3724_1), .IN4(~na1153_1), .IN5(1'b1), .IN6(na1136_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y104     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1153_1 ( .OUT(na1153_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2458_2), .IN6(1'b0), .IN7(~na2426_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x140y105     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_1 ( .OUT(na1154_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1155_1), .IN6(na3729_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y99     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_1 ( .OUT(na1155_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2459_1), .IN6(1'b0), .IN7(~na2427_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x136y98     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1156_1 ( .OUT(na1156_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3730_1), .IN6(~na1157_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x121y92     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_1 ( .OUT(na1157_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2460_2), .IN4(~na2428_2), .IN5(1'b1), .IN6(~na2416_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y102     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1158_1 ( .OUT(na1158_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1159_1), .IN8(na3733_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x110y103     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1159_1 ( .OUT(na1159_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2461_1), .IN4(~na2429_1), .IN5(1'b1), .IN6(~na2416_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x136y95     80'h00_0018_00_0040_0A51_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1160_1 ( .OUT(na1160_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4258_2), .IN5(~na1161_1), .IN6(1'b0), .IN7(na3734_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y91     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_1 ( .OUT(na1161_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2462_2), .IN6(1'b0), .IN7(~na2430_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y92     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1162_1 ( .OUT(na1162_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1163_1), .IN6(na3735_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y83     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_1 ( .OUT(na1163_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4327_2), .IN8(~na2431_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x131y98     80'h00_0018_00_0040_0C13_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1164_1 ( .OUT(na1164_1), .IN1(~na1165_1), .IN2(na3736_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1136_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y95     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2432_1), .IN6(~na2464_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x130y90     80'h00_0018_00_0040_0C4C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1166_1 ( .OUT(na1166_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1167_1), .IN4(na3737_1), .IN5(1'b1), .IN6(~na1136_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y79     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1167_1 ( .OUT(na1167_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4310_2), .IN5(~na4317_2), .IN6(1'b0), .IN7(~na2465_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x139y99     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3762_2), .IN8(~na1169_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y102     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1169_1 ( .OUT(na1169_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na2434_1), .IN7(1'b0), .IN8(~na2466_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x137y96     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_1 ( .OUT(na1170_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3767_2), .IN8(~na1171_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x136y100     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_1 ( .OUT(na1171_1), .IN1(~na2435_1), .IN2(~na2467_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2416_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x138y97     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1172_1 ( .OUT(na1172_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3768_1), .IN8(~na1173_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x126y100     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_1 ( .OUT(na1173_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4330_2), .IN4(~na2436_1), .IN5(1'b1), .IN6(~na2416_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y99     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1174_1 ( .OUT(na1174_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1175_1), .IN8(na3771_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y101     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1175_1 ( .OUT(na1175_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2437_1), .IN6(~na2469_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y93     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1176_1 ( .OUT(na1176_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3772_1), .IN8(~na1177_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y90     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1177_1 ( .OUT(na1177_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na4318_2), .IN7(1'b0), .IN8(~na2470_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x132y83     80'h00_0018_00_0040_0C4C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1178_1 ( .OUT(na1178_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1179_1), .IN4(na3773_2), .IN5(1'b1), .IN6(~na1136_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y77     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1179_1 ( .OUT(na1179_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2439_2), .IN6(~na2471_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x136y92     80'h00_0018_00_0040_0C8C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1180_1 ( .OUT(na1180_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3774_2), .IN4(~na1181_1), .IN5(1'b1), .IN6(na1136_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y94     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1181_1 ( .OUT(na1181_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na4332_2), .IN6(1'b0), .IN7(~na2440_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y88     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1182_1 ( .OUT(na1182_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1183_1), .IN6(na3775_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x113y81     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1183_1 ( .OUT(na1183_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2473_1), .IN6(1'b0), .IN7(~na2441_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y107     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1184_1 ( .OUT(na1184_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1185_1), .IN6(na3801_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x119y105     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1185_1 ( .OUT(na1185_1), .IN1(~na2474_1), .IN2(~na2442_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2416_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y103     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1186_1 ( .OUT(na1186_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3806_1), .IN8(~na1187_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x132y100     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1187_1 ( .OUT(na1187_1), .IN1(~na2443_1), .IN2(~na4333_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2416_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x133y103     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1188_1 ( .OUT(na1188_1), .IN1(1'b1), .IN2(~na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1189_1), .IN6(na3807_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y107     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1189_1 ( .OUT(na1189_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4310_2), .IN5(~na2444_2), .IN6(1'b0), .IN7(~na2476_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y103     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1190_1 ( .OUT(na1190_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3810_1), .IN8(~na1191_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y110     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1191_1 ( .OUT(na1191_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2445_1), .IN6(~na4334_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x134y102     80'h00_0018_00_0040_0C13_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1192_1 ( .OUT(na1192_1), .IN1(~na1193_1), .IN2(na3811_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1136_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y93     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1193_1 ( .OUT(na1193_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2478_1), .IN6(~na2446_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x126y97     80'h00_0018_00_0040_0C8C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1194_1 ( .OUT(na1194_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3812_1), .IN4(~na1195_1), .IN5(1'b1), .IN6(na1136_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y86     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1195_1 ( .OUT(na1195_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(~na2479_2), .IN7(1'b0), .IN8(~na2447_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y97     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1196_1 ( .OUT(na1196_1), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3813_2), .IN8(~na1197_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y94     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1197_1 ( .OUT(na1197_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2480_1), .IN6(1'b0), .IN7(~na2448_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y98     80'h00_0018_00_0040_0A51_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1198_1 ( .OUT(na1198_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4258_2), .IN5(~na1199_1), .IN6(1'b0), .IN7(na3814_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x107y91     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_1 ( .OUT(na1199_1), .IN1(~na2481_1), .IN2(~na4320_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2416_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y72     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1200_1 ( .OUT(na1200_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na539_2), .IN7(1'b1), .IN8(na1900_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y72     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1201_4 ( .OUT(na1201_2), .IN1(1'b1), .IN2(~na539_2), .IN3(1'b1), .IN4(na1900_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y72     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1202_1 ( .OUT(na1202_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3235_2), .IN6(~na539_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x145y94     80'h00_0018_00_0000_0EEE_DC53
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1203_1 ( .OUT(na1203_1), .IN1(1'b0), .IN2(~na3944_1), .IN3(~na3959_2), .IN4(1'b0), .IN5(1'b0), .IN6(na3962_1), .IN7(~na3959_1),
                      .IN8(na3960_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x149y73     80'h00_0060_00_0000_0C08_FF2A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1206_4 ( .OUT(na1206_2), .IN1(na1207_2), .IN2(1'b1), .IN3(na1930_1), .IN4(~na1932_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y77     80'h00_0060_00_0000_0C08_FF13
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1207_4 ( .OUT(na1207_2), .IN1(1'b1), .IN2(~na1929_1), .IN3(~na1930_2), .IN4(~na1932_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y83     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1208_1 ( .OUT(na1208_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1209_1), .IN6(1'b1), .IN7(na1930_1), .IN8(na1932_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y83     80'h00_0018_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1209_1 ( .OUT(na1209_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1929_1), .IN7(na1930_2), .IN8(~na1932_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y77     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1211_4 ( .OUT(na1211_2), .IN1(na1207_2), .IN2(1'b1), .IN3(na538_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y79     80'h00_0018_00_0000_0C88_4AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1212_1 ( .OUT(na1212_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1213_2), .IN6(1'b1), .IN7(~na1930_1), .IN8(na1932_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y79     80'h00_0060_00_0000_0C08_FF23
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1213_4 ( .OUT(na1213_2), .IN1(1'b1), .IN2(~na1929_1), .IN3(na1930_2), .IN4(~na1932_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x147y96     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1214_1 ( .OUT(na1214_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3950_1), .IN6(na3281_1), .IN7(1'b0), .IN8(na1932_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y89     80'h00_0018_00_0000_0888_8811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1217_1 ( .OUT(na1217_1), .IN1(~na3952_1), .IN2(~na3954_2), .IN3(~na3956_2), .IN4(~na3958_1), .IN5(na3955_1), .IN6(na3953_2),
                      .IN7(na3957_1), .IN8(na3951_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y75     80'h00_0060_00_0000_0C08_FF4A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1219_4 ( .OUT(na1219_2), .IN1(na1207_2), .IN2(1'b1), .IN3(~na1930_1), .IN4(na1932_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y77     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1220_1 ( .OUT(na1220_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1213_2), .IN6(1'b1), .IN7(na538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y77     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1222_4 ( .OUT(na1222_2), .IN1(1'b1), .IN2(na1223_1), .IN3(na538_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y80     80'h00_0018_00_0000_0C88_1CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1223_1 ( .OUT(na1223_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1929_1), .IN7(~na1930_2), .IN8(~na1932_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y83     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1224_4 ( .OUT(na1224_2), .IN1(na1209_1), .IN2(1'b1), .IN3(na538_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y74     80'h00_0060_00_0000_0C08_FF2C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1226_4 ( .OUT(na1226_2), .IN1(1'b1), .IN2(na1223_1), .IN3(na1930_1), .IN4(~na1932_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y82     80'h00_0018_00_0000_0C88_2AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1227_1 ( .OUT(na1227_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1209_1), .IN6(1'b1), .IN7(na1930_1), .IN8(~na1932_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y82     80'h00_0060_00_0000_0C08_FF4A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1229_4 ( .OUT(na1229_2), .IN1(na1209_1), .IN2(1'b1), .IN3(~na1930_1), .IN4(na1932_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y82     80'h00_0060_00_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1230_4 ( .OUT(na1230_2), .IN1(na1207_2), .IN2(1'b1), .IN3(na1930_1), .IN4(na1932_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y85     80'h00_0018_00_0000_0C88_4CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1232_1 ( .OUT(na1232_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1223_1), .IN7(~na1930_1), .IN8(na1932_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y80     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1233_4 ( .OUT(na1233_2), .IN1(1'b1), .IN2(na1223_1), .IN3(na1930_1), .IN4(na1932_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y85     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1235_1 ( .OUT(na1235_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1213_2), .IN6(1'b1), .IN7(na1930_1), .IN8(na1932_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y78     80'h00_0060_00_0000_0C08_FF2A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1236_4 ( .OUT(na1236_2), .IN1(na1213_2), .IN2(1'b1), .IN3(na1930_1), .IN4(~na1932_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x145y93     80'h00_0018_00_0000_0EEE_DA55
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1237_1 ( .OUT(na1237_1), .IN1(~na3963_1), .IN2(1'b0), .IN3(~na3975_2), .IN4(1'b0), .IN5(na3978_2), .IN6(1'b0), .IN7(~na3975_1),
                      .IN8(na3976_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y93     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_1 ( .OUT(na1239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3091_1), .IN8(na1230_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x142y88     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1242_4 ( .OUT(na1242_2), .IN1(~na1206_2), .IN2(~na2407_1), .IN3(~na1224_2), .IN4(~na3059_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x143y87     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1243_1 ( .OUT(na1243_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1219_2), .IN6(~na2899_1), .IN7(~na1212_1),
                      .IN8(~na2995_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x144y89     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1244_1 ( .OUT(na1244_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1232_1), .IN6(~na3067_1), .IN7(~na1220_1),
                      .IN8(~na3003_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x144y92     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1245_4 ( .OUT(na1245_2), .IN1(~na2939_1), .IN2(~na1229_2), .IN3(~na3083_2), .IN4(~na1233_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x144y84     80'h00_0018_00_0000_0EEE_5E55
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1248_1 ( .OUT(na1248_1), .IN1(~na3979_1), .IN2(1'b0), .IN3(~na3990_2), .IN4(1'b0), .IN5(na3993_1), .IN6(na3991_1), .IN7(~na3990_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x143y76     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1251_4 ( .OUT(na1251_2), .IN1(na2900_2), .IN2(1'b1), .IN3(na4261_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x146y80     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1254_1 ( .OUT(na1254_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2988_2), .IN6(~na1226_2), .IN7(~na1212_1),
                      .IN8(~na2996_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x141y81     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1255_1 ( .OUT(na1255_1), .IN1(~na3052_2), .IN2(~na1227_1), .IN3(~na3092_2), .IN4(~na1230_2), .IN5(~na2980_2), .IN6(~na4267_2),
                      .IN7(~na1235_1), .IN8(~na4295_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x145y92     80'h00_0018_00_0000_0EEE_C55D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1260_1 ( .OUT(na1260_1), .IN1(~na4006_2), .IN2(na4009_1), .IN3(~na3994_1), .IN4(1'b0), .IN5(~na4006_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na4007_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y86     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1262_4 ( .OUT(na1262_2), .IN1(na2901_1), .IN2(1'b1), .IN3(na4261_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x141y86     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1265_4 ( .OUT(na1265_2), .IN1(~na3005_1), .IN2(~na4262_2), .IN3(~na3093_1), .IN4(~na1230_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x143y83     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1266_1 ( .OUT(na1266_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1211_2), .IN6(~na4379_2), .IN7(~na2981_1),
                      .IN8(~na1236_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x142y88     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1267_1 ( .OUT(na1267_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3053_1), .IN6(~na1227_1), .IN7(~na1235_1),
                      .IN8(~na1923_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x145y84     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1268_4 ( .OUT(na1268_2), .IN1(~na2989_1), .IN2(~na1226_2), .IN3(~na1208_1), .IN4(~na3077_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y76     80'h00_0018_00_0000_0888_8812
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_1 ( .OUT(na1271_1), .IN1(na1277_1), .IN2(~na4011_1), .IN3(~na4013_1), .IN4(~na4015_2), .IN5(na4012_1), .IN6(na4010_1),
                      .IN7(na4014_1), .IN8(na1276_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x142y72     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1276_1 ( .OUT(na1276_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4263_2), .IN6(~na3046_2), .IN7(~na1220_1),
                      .IN8(~na3006_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y75     80'h00_0018_00_0000_0888_8811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1277_1 ( .OUT(na1277_1), .IN1(~na4021_2), .IN2(~na4025_2), .IN3(~na4023_2), .IN4(~na4019_2), .IN5(na4018_1), .IN6(na4020_1),
                      .IN7(na4024_1), .IN8(na4022_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y74     80'h00_0018_00_0000_0888_8821
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1282_1 ( .OUT(na1282_1), .IN1(~na4029_2), .IN2(~na4027_2), .IN3(na1288_1), .IN4(~na4031_2), .IN5(na1287_1), .IN6(na4026_1),
                      .IN7(na4028_1), .IN8(na4030_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x145y73     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1287_1 ( .OUT(na1287_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2943_1), .IN6(~na1229_2), .IN7(~na2983_1),
                      .IN8(~na1236_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y71     80'h00_0018_00_0000_0888_8811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1288_1 ( .OUT(na1288_1), .IN1(~na4035_2), .IN2(~na4039_1), .IN3(~na4037_1), .IN4(~na4041_1), .IN5(na4034_1), .IN6(na4036_2),
                      .IN7(na4040_2), .IN8(na4038_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x145y83     80'h00_0018_00_0000_0EEE_5A5D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1293_1 ( .OUT(na1293_1), .IN1(~na4042_1), .IN2(na4057_2), .IN3(~na4054_2), .IN4(1'b0), .IN5(na4055_1), .IN6(1'b0), .IN7(~na4054_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y73     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1295_1 ( .OUT(na1295_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1206_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2412_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x139y76     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1298_4 ( .OUT(na1298_2), .IN1(~na1232_1), .IN2(~na3072_2), .IN3(~na4261_2), .IN4(~na2904_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x145y77     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1299_1 ( .OUT(na1299_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3088_2), .IN6(~na4266_2), .IN7(~na1212_1),
                      .IN8(~na4354_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x145y80     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1300_4 ( .OUT(na1300_2), .IN1(~na3008_2), .IN2(~na4262_2), .IN3(~na1208_1), .IN4(~na3080_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x142y82     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1301_4 ( .OUT(na1301_2), .IN1(~na2944_2), .IN2(~na1229_2), .IN3(~na3096_2), .IN4(~na1230_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x146y76     80'h00_0018_00_0000_0EEE_DBED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1304_1 ( .OUT(na1304_1), .IN1(~na4058_1), .IN2(na1312_2), .IN3(na4415_2), .IN4(na1313_1), .IN5(na4068_2), .IN6(~na1316_1),
                      .IN7(~na4067_2), .IN8(na4066_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x141y72     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1306_4 ( .OUT(na1306_2), .IN1(na3089_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1233_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y75     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1309_1 ( .OUT(na1309_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1212_1), .IN8(na3001_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y72     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1312_4 ( .OUT(na1312_2), .IN1(na1206_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2413_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y82     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3065_1), .IN7(na1224_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x141y74     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1316_1 ( .OUT(na1316_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1219_2), .IN6(~na4346_2), .IN7(~na4353_2),
                      .IN8(~na1236_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y68     80'h00_0018_00_0040_0C65_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1317_1 ( .OUT(na1317_1), .IN1(na4071_1), .IN2(1'b1), .IN3(~na3151_1), .IN4(1'b0), .IN5(~na4382_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3150_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x129y66     80'h00_0018_00_0040_0C9D_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1318_1 ( .OUT(na1318_1), .IN1(~na4072_2), .IN2(1'b0), .IN3(na3151_2), .IN4(~na4383_2), .IN5(~na4381_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3150_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x135y75     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1319_1 ( .OUT(na1319_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1126_2), .IN7(1'b1), .IN8(~na4310_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x127y70     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1320_4 ( .OUT(na1320_2), .IN1(1'b1), .IN2(~na1126_2), .IN3(1'b1), .IN4(na1871_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x129y74     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1321_1 ( .OUT(na1321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1126_2), .IN7(1'b1), .IN8(na1871_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y69     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1322_4 ( .OUT(na1322_2), .IN1(1'b1), .IN2(~na1126_2), .IN3(na1873_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y81     80'h00_0018_00_0000_0888_AC84
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_1 ( .OUT(na1323_1), .IN1(~na4388_2), .IN2(na1325_1), .IN3(na3170_2), .IN4(na3172_2), .IN5(1'b1), .IN6(na3185_1), .IN7(na3170_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y68     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1324_4 ( .OUT(na1324_2), .IN1(na4384_2), .IN2(na1325_1), .IN3(na3170_2), .IN4(na3172_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y72     80'h00_0018_00_0000_0888_8218
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_1 ( .OUT(na1325_1), .IN1(na3175_1), .IN2(na1328_2), .IN3(~na4387_2), .IN4(~na3182_1), .IN5(na3175_2), .IN6(~na3181_2),
                      .IN7(na3174_2), .IN8(na3182_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y66     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1328_4 ( .OUT(na1328_2), .IN1(~na3178_1), .IN2(~na3176_1), .IN3(~na3180_1), .IN4(~na3173_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y66     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1329_1 ( .OUT(na1329_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4073_2), .IN7(~na3170_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y66     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1330_4 ( .OUT(na1330_2), .IN1(na1886_1), .IN2(~na4073_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y66     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1331_1 ( .OUT(na1331_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1886_2), .IN6(~na4073_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y67     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1332_4 ( .OUT(na1332_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1333_1), .IN4(~na3173_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y69     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1), .IN1(1'b1), .IN2(na3185_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na4076_2), .IN6(na1325_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y70     80'h00_0018_00_0000_0888_2121
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1334_1 ( .OUT(na1334_1), .IN1(~na3175_1), .IN2(~na3181_1), .IN3(na1336_2), .IN4(~na3182_1), .IN5(~na3175_2), .IN6(~na3181_2),
                      .IN7(na3174_2), .IN8(~na3182_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y67     80'h00_0060_00_0000_0C08_FF48
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1336_4 ( .OUT(na1336_2), .IN1(na3178_1), .IN2(na3176_1), .IN3(~na3180_1), .IN4(na3173_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y68     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1337_1 ( .OUT(na1337_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1876_1), .IN7(~na1333_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y69     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1338_4 ( .OUT(na1338_2), .IN1(1'b1), .IN2(na1876_2), .IN3(~na1333_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y67     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1339_1 ( .OUT(na1339_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1878_1), .IN6(1'b1), .IN7(~na1333_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y69     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1340_1 ( .OUT(na1340_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1878_2), .IN6(1'b1), .IN7(~na1333_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y71     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1341_1 ( .OUT(na1341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1880_1), .IN7(~na1333_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y72     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1342_4 ( .OUT(na1342_2), .IN1(1'b1), .IN2(na1880_2), .IN3(~na1333_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y72     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1343_1 ( .OUT(na1343_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1882_1), .IN6(1'b1), .IN7(~na1333_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y76     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1344_4 ( .OUT(na1344_2), .IN1(na1882_2), .IN2(1'b1), .IN3(~na1333_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y73     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1884_1), .IN7(~na1333_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y74     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1346_4 ( .OUT(na1346_2), .IN1(1'b1), .IN2(na1884_2), .IN3(~na1333_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y76     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1347_1 ( .OUT(na1347_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3185_1), .IN7(na3184_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x147y67     80'h00_0018_00_0040_0C68_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1348_1 ( .OUT(na1348_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na2399_1), .IN5(1'b1), .IN6(~na4391_2), .IN7(na3223_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y88     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1349_1 ( .OUT(na1349_1), .IN1(1'b1), .IN2(na539_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2400_2), .IN6(na1941_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y89     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1350_1 ( .OUT(na1350_1), .IN1(1'b1), .IN2(na539_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2401_2), .IN8(na1946_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x146y94     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_1 ( .OUT(na1351_1), .IN1(1'b1), .IN2(na539_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2402_2), .IN6(na1941_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y94     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1352_1 ( .OUT(na1352_1), .IN1(1'b1), .IN2(~na539_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1943_2), .IN8(na2403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y91     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_1 ( .OUT(na1353_1), .IN1(1'b1), .IN2(~na539_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1943_1), .IN8(na2404_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y90     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1354_1 ( .OUT(na1354_1), .IN1(1'b1), .IN2(~na539_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1945_2), .IN6(na2405_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x146y92     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1355_1 ( .OUT(na1355_1), .IN1(1'b1), .IN2(~na539_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1945_1), .IN6(na1911_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y65     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1356_4 ( .OUT(na1356_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na3212_2), .IN4(~na4271_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x146y67     80'h00_0018_00_0040_0C76_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1357_1 ( .OUT(na1357_1), .IN1(1'b1), .IN2(~na4392_2), .IN3(~na3223_2), .IN4(1'b0), .IN5(~na1358_1), .IN6(1'b1), .IN7(na3223_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y67     80'h00_0018_00_0000_0888_1828
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1358_1 ( .OUT(na1358_1), .IN1(na3214_1), .IN2(na1361_1), .IN3(na3216_1), .IN4(~na3220_1), .IN5(na3214_2), .IN6(na3213_1),
                      .IN7(~na3216_2), .IN8(~na3220_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y66     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1361_1 ( .OUT(na1361_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3215_2), .IN6(~na3217_1), .IN7(~na3212_2),
                      .IN8(~na3219_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y65     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1362_1 ( .OUT(na1362_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1890_1), .IN6(1'b1), .IN7(~na1357_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y66     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1363_4 ( .OUT(na1363_2), .IN1(na1890_2), .IN2(1'b1), .IN3(~na1357_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x140y68     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1892_1), .IN7(~na1357_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y66     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1365_4 ( .OUT(na1365_2), .IN1(1'b1), .IN2(na1892_2), .IN3(~na1357_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y68     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_1 ( .OUT(na1366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1894_1), .IN6(1'b1), .IN7(~na1357_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y67     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1367_4 ( .OUT(na1367_2), .IN1(na1894_2), .IN2(1'b1), .IN3(~na1357_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y69     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1368_1 ( .OUT(na1368_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1896_1), .IN7(~na1357_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y66     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1369_4 ( .OUT(na1369_2), .IN1(1'b1), .IN2(na1896_2), .IN3(~na1357_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y71     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1370_1 ( .OUT(na1370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1898_1), .IN6(1'b1), .IN7(~na1357_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x143y68     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1371_4 ( .OUT(na1371_2), .IN1(na1898_2), .IN2(1'b1), .IN3(~na1357_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x147y66     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1372_1 ( .OUT(na1372_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na4391_2), .IN7(na3223_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x103y85     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1373_4 ( .OUT(na1373_2), .IN1(~na4304_2), .IN2(~na1957_2), .IN3(na3169_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y69     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1374_1 ( .OUT(na1374_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1957_2), .IN7(na1958_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y98     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1375_1 ( .OUT(na1375_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1377_2), .IN6(~na1937_2), .IN7(na4274_2),
                      .IN8(~na4297_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y102     80'h00_0018_00_0000_0C88_32FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1376_1 ( .OUT(na1376_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1373_2), .IN6(~na1937_1), .IN7(1'b1), .IN8(~na1938_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y95     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1377_4 ( .OUT(na1377_2), .IN1(~na1935_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y68     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1378_1 ( .OUT(na1378_1), .IN1(1'b1), .IN2(na539_2), .IN3(1'b1), .IN4(na1379_2), .IN5(na1358_1), .IN6(na4302_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y70     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1379_4 ( .OUT(na1379_2), .IN1(~na1380_1), .IN2(~na4391_2), .IN3(na3223_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y69     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1380_1 ( .OUT(na1380_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3235_1), .IN6(na3234_1), .IN7(1'b1), .IN8(na4394_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y87     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1381_1 ( .OUT(na1381_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4389_2), .IN6(na1325_1), .IN7(~na3184_2),
                      .IN8(na3277_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y87     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1382_4 ( .OUT(na1382_2), .IN1(1'b1), .IN2(na1383_1), .IN3(1'b1), .IN4(~na3695_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x147y70     80'h00_0018_00_0000_0888_DFA3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1383_1 ( .OUT(na1383_1), .IN1(1'b0), .IN2(~na4391_2), .IN3(na3277_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(~na3223_2),
                      .IN8(na4272_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y73     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1384_1 ( .OUT(na1384_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1385_1), .IN8(na4079_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x90y75     80'h00_0018_00_0040_0CCB_5300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1385_1 ( .OUT(na1385_1), .IN1(na4390_2), .IN2(na1334_1), .IN3(1'b1), .IN4(~na3211_2), .IN5(1'b1), .IN6(~na3185_1), .IN7(~na3184_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y89     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1386_4 ( .OUT(na1386_2), .IN1(1'b1), .IN2(na1387_1), .IN3(na1389_1), .IN4(na1388_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y98     80'h00_0018_00_0000_0C88_C2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1373_2), .IN6(~na1937_1), .IN7(1'b1), .IN8(na1938_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y98     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1388_4 ( .OUT(na1388_2), .IN1(na1935_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y97     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1389_1 ( .OUT(na1389_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1935_1), .IN6(na1937_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y91     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1390_4 ( .OUT(na1390_2), .IN1(na1377_2), .IN2(na1387_1), .IN3(na1389_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y94     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1391_1 ( .OUT(na1391_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1387_1), .IN7(na1389_1), .IN8(na1392_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y98     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1392_4 ( .OUT(na1392_2), .IN1(na1935_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y95     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1393_4 ( .OUT(na1393_2), .IN1(~na1935_2), .IN2(na1387_1), .IN3(na1389_1), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y94     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1394_1 ( .OUT(na1394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1387_1), .IN7(na1395_1), .IN8(na1388_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y99     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1395_1 ( .OUT(na1395_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_1), .IN6(na1937_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y91     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1396_1 ( .OUT(na1396_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1377_2), .IN6(na1387_1), .IN7(na1395_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y90     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1397_4 ( .OUT(na1397_2), .IN1(1'b1), .IN2(na1387_1), .IN3(na1395_1), .IN4(na1392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y94     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1398_4 ( .OUT(na1398_2), .IN1(~na1935_2), .IN2(na1387_1), .IN3(na1395_1), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y95     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1399_1 ( .OUT(na1399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1387_1), .IN7(na1400_2), .IN8(na1388_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y97     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1400_4 ( .OUT(na1400_2), .IN1(na1935_1), .IN2(~na1937_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y91     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1401_4 ( .OUT(na1401_2), .IN1(na1377_2), .IN2(na1387_1), .IN3(na1400_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y93     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1402_1 ( .OUT(na1402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1387_1), .IN7(na1400_2), .IN8(na1392_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y89     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1403_4 ( .OUT(na1403_2), .IN1(~na1935_2), .IN2(na1387_1), .IN3(na1400_2), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y96     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1404_1 ( .OUT(na1404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_1), .IN6(~na1937_2), .IN7(na4276_2),
                      .IN8(na1388_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y99     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1405_4 ( .OUT(na1405_2), .IN1(1'b1), .IN2(na1406_1), .IN3(na1395_1), .IN4(na1388_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y100     80'h00_0018_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1406_1 ( .OUT(na1406_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1373_2), .IN6(na1937_1), .IN7(1'b1), .IN8(~na1938_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y93     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1407_4 ( .OUT(na1407_2), .IN1(~na1935_2), .IN2(na1406_1), .IN3(na1389_1), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y96     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1408_4 ( .OUT(na1408_2), .IN1(1'b1), .IN2(na1406_1), .IN3(na1389_1), .IN4(na1392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y95     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1409_1 ( .OUT(na1409_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1377_2), .IN6(na1406_1), .IN7(na1389_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y84     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1410_4 ( .OUT(na1410_2), .IN1(1'b1), .IN2(na535_2), .IN3(na4275_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y94     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_1 ( .OUT(na1411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_1), .IN6(~na1937_2), .IN7(na4276_2),
                      .IN8(na1392_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y93     80'h00_0060_00_0000_0C08_FF22
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1412_4 ( .OUT(na1412_2), .IN1(na1377_2), .IN2(~na1937_2), .IN3(na4276_2), .IN4(~na4297_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y94     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1413_4 ( .OUT(na1413_2), .IN1(na1377_2), .IN2(na1406_1), .IN3(na1395_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y98     80'h00_0018_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1414_1 ( .OUT(na1414_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_2), .IN6(na1406_1), .IN7(na1400_2),
                      .IN8(~na1934_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y99     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1415_1 ( .OUT(na1415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1406_1), .IN7(na1400_2), .IN8(na1392_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y95     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1416_4 ( .OUT(na1416_2), .IN1(na1377_2), .IN2(na1406_1), .IN3(na1400_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y103     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1417_1 ( .OUT(na1417_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1406_1), .IN7(na1400_2), .IN8(na1388_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y95     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1418_4 ( .OUT(na1418_2), .IN1(~na1935_2), .IN2(na1406_1), .IN3(na1395_1), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y98     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1419_4 ( .OUT(na1419_2), .IN1(1'b1), .IN2(na1406_1), .IN3(na1395_1), .IN4(na1392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y104     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1420_1 ( .OUT(na1420_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_1), .IN6(~na1937_2), .IN7(na4278_2),
                      .IN8(na1388_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y98     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1421_1 ( .OUT(na1421_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1376_1), .IN7(na1389_1), .IN8(na1392_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y94     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1422_4 ( .OUT(na1422_2), .IN1(na1377_2), .IN2(na1376_1), .IN3(na1389_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y99     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1423_4 ( .OUT(na1423_2), .IN1(1'b1), .IN2(na1376_1), .IN3(na1389_1), .IN4(na1388_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y94     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1424_4 ( .OUT(na1424_2), .IN1(1'b1), .IN2(na535_2), .IN3(1'b1), .IN4(na4277_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y99     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1425_4 ( .OUT(na1425_2), .IN1(~na1935_1), .IN2(~na1937_2), .IN3(na4278_2), .IN4(na1392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y98     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1426_1 ( .OUT(na1426_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1377_2), .IN6(~na1937_2), .IN7(na4278_2),
                      .IN8(~na4297_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y98     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1427_4 ( .OUT(na1427_2), .IN1(~na1935_2), .IN2(na1376_1), .IN3(na1389_1), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y96     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1428_4 ( .OUT(na1428_2), .IN1(na1377_2), .IN2(na1376_1), .IN3(na1400_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y101     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1429_1 ( .OUT(na1429_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1376_1), .IN7(na1400_2), .IN8(na1388_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y97     80'h00_0018_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1430_1 ( .OUT(na1430_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_2), .IN6(na1376_1), .IN7(na1395_1),
                      .IN8(~na1934_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y96     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1431_4 ( .OUT(na1431_2), .IN1(1'b1), .IN2(na1376_1), .IN3(na1395_1), .IN4(na1392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y97     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1432_1 ( .OUT(na1432_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1377_2), .IN6(na1376_1), .IN7(na1395_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y99     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1433_4 ( .OUT(na1433_2), .IN1(1'b1), .IN2(na1376_1), .IN3(na1395_1), .IN4(na1388_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y99     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1434_1 ( .OUT(na1434_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1376_1), .IN7(na1400_2), .IN8(na1392_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x89y71     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1435_4 ( .OUT(na1435_2), .IN1(na4270_2), .IN2(~na3185_1), .IN3(~na3184_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y68     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1436_1 ( .OUT(na1436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3185_1), .IN7(na3184_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y84     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1437_4 ( .OUT(na1437_2), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x131y84     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1438_4 ( .OUT(na1438_2), .IN1(1'b1), .IN2(~na543_2), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y80     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1439_4 ( .OUT(na1439_2), .IN1(1'b1), .IN2(1'b1), .IN3(na17_1), .IN4(na4082_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x140y76     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1440_1 ( .OUT(na1440_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na21_2), .IN6(~na1126_2), .IN7(1'b0), .IN8(~na1441_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y108     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1441_4 ( .OUT(na1441_2), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x137y81     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1442_4 ( .OUT(na1442_2), .IN1(~na4255_2), .IN2(~na16_2), .IN3(1'b0), .IN4(~na1441_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x139y75     80'h00_0018_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1443_1 ( .OUT(na1443_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na21_2), .IN6(na4268_2), .IN7(na4085_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x138y81     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1445_1 ( .OUT(na1445_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na4083_1), .IN6(na2416_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x132y79     80'h00_0018_00_0040_0C27_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1446_1 ( .OUT(na1446_1), .IN1(na4255_2), .IN2(~na543_2), .IN3(na4088_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na16_2), .IN7(1'b1),
                      .IN8(~na4310_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x139y70     80'h00_0060_00_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1447_4 ( .OUT(na1447_2), .IN1(na1319_1), .IN2(~na16_2), .IN3(na4089_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x138y77     80'h00_0018_00_0040_0C06_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1449_1 ( .OUT(na1449_1), .IN1(1'b0), .IN2(na1126_2), .IN3(na4269_2), .IN4(1'b0), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(na19_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x136y84     80'h00_0018_00_0000_0888_FE53
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1450_1 ( .OUT(na1450_1), .IN1(1'b0), .IN2(~na1437_2), .IN3(~na26_2), .IN4(1'b0), .IN5(na4170_2), .IN6(na543_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y84     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(1'b0), .IN6(na1126_2), .IN7(1'b0), .IN8(na1441_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x137y78     80'h00_0018_00_0000_0C88_CBFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1452_1 ( .OUT(na1452_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1319_1), .IN6(~na16_2), .IN7(1'b0), .IN8(na1453_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x132y68     80'h00_0018_00_0040_0C05_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1453_1 ( .OUT(na1453_1), .IN1(na4093_1), .IN2(1'b0), .IN3(na3151_1), .IN4(1'b0), .IN5(na4382_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na3150_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y103     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1454_1 ( .OUT(na1454_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na534_2), .IN7(~na3169_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x144y71     80'h00_0060_00_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1455_4 ( .OUT(na1455_2), .IN1(na537_1), .IN2(~na1957_2), .IN3(na1958_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x132y81     80'h00_0018_00_0040_0C2E_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1456_1 ( .OUT(na1456_1), .IN1(1'b0), .IN2(~na543_2), .IN3(na4088_2), .IN4(na4256_2), .IN5(1'b1), .IN6(na2416_2), .IN7(1'b1),
                      .IN8(~na19_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x129y68     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1457_1 ( .OUT(na1457_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1386_2), .IN6(1'b0), .IN7(na1958_1), .IN8(~na4303_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x127y77     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1458_4 ( .OUT(na1458_2), .IN1(1'b1), .IN2(~na543_2), .IN3(~na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x135y80     80'h00_0018_00_0000_0888_FEAE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1459_1 ( .OUT(na1459_1), .IN1(na21_2), .IN2(na4268_2), .IN3(na17_1), .IN4(1'b0), .IN5(na4380_2), .IN6(na1126_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x104y98     80'h00_0018_00_0000_0888_FD55
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1460_1 ( .OUT(na1460_1), .IN1(~na1458_2), .IN2(1'b0), .IN3(~na26_2), .IN4(1'b0), .IN5(~na4257_2), .IN6(na57_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y98     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1461_4 ( .OUT(na1461_2), .IN1(1'b1), .IN2(na1406_1), .IN3(na1389_1), .IN4(na1388_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x105y97     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1462_1 ( .OUT(na1462_1), .IN1(na4100_2), .IN2(na543_2), .IN3(~na26_2), .IN4(1'b0), .IN5(~na4257_2), .IN6(na57_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y95     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1464_4 ( .OUT(na1464_2), .IN1(~na1935_2), .IN2(na1376_1), .IN3(na1400_2), .IN4(~na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y102     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1465_1 ( .OUT(na1465_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1935_1), .IN6(~na1937_2), .IN7(na4274_2),
                      .IN8(na1388_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y95     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1466_4 ( .OUT(na1466_2), .IN1(1'b1), .IN2(na535_2), .IN3(1'b1), .IN4(na4273_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y98     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1467_4 ( .OUT(na1467_2), .IN1(~na1935_1), .IN2(~na1937_2), .IN3(na4274_2), .IN4(na1392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x121y68     80'h00_0018_00_0040_0C03_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1468_1 ( .OUT(na1468_1), .IN1(na4101_1), .IN2(na4102_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3132_2), .IN7(na3130_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x99y115     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1469_1 ( .OUT(na1469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na959_1), .IN6(na3202_2), .IN7(na2762_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y110     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1470_1 ( .OUT(na1470_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2763_1), .IN7(na3203_1), .IN8(na1003_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y115     80'h00_0018_00_0000_0666_AC9C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1471_1 ( .OUT(na1471_1), .IN1(1'b0), .IN2(na1014_2), .IN3(~na1016_1), .IN4(na1013_2), .IN5(1'b0), .IN6(na3204_2), .IN7(na2764_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y116     80'h00_0018_00_0000_0666_AC9C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1473_1 ( .OUT(na1473_1), .IN1(1'b0), .IN2(na1020_1), .IN3(na2765_1), .IN4(~na996_2), .IN5(1'b0), .IN6(na3205_1), .IN7(na1016_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x100y115     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1475_4 ( .OUT(na1475_2), .IN1(na1026_2), .IN2(~na2766_2), .IN3(na1016_1), .IN4(~na3206_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x89y104     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1476_1 ( .OUT(na1476_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3207_1), .IN6(~na2767_1), .IN7(na1030_1),
                      .IN8(na4253_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x102y107     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1477_1 ( .OUT(na1477_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3208_2), .IN6(na2768_2), .IN7(1'b0), .IN8(na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x89y107     80'h00_0018_00_0000_0666_A59C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1478_1 ( .OUT(na1478_1), .IN1(1'b0), .IN2(na1035_1), .IN3(na1030_1), .IN4(~na1015_1), .IN5(~na2769_1), .IN6(1'b0), .IN7(na3209_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x89y109     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1480_1 ( .OUT(na1480_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2738_2), .IN7(na215_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x94y99     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1481_4 ( .OUT(na1481_2), .IN1(1'b0), .IN2(na2739_1), .IN3(1'b0), .IN4(na263_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x100y82     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1482_1 ( .OUT(na1482_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2740_1), .IN7(1'b0), .IN8(na275_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x89y115     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1483_4 ( .OUT(na1483_2), .IN1(na2741_1), .IN2(1'b0), .IN3(na281_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y79     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1484_1 ( .OUT(na1484_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2742_2), .IN6(1'b0), .IN7(na293_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y85     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1485_1 ( .OUT(na1485_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na298_1), .IN8(na2743_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x97y90     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1486_1 ( .OUT(na1486_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(1'b0), .IN7(1'b0), .IN8(na2424_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x100y70     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1487_4 ( .OUT(na1487_2), .IN1(na312_1), .IN2(1'b0), .IN3(na2745_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x128y110     80'h00_0060_00_0000_0C06_FF9A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1488_4 ( .OUT(na1488_2), .IN1(na808_2), .IN2(1'b0), .IN3(na848_1), .IN4(~na2746_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y106     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1489_4 ( .OUT(na1489_2), .IN1(na852_1), .IN2(1'b0), .IN3(na2427_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x142y110     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1490_4 ( .OUT(na1490_2), .IN1(na808_2), .IN2(~na2748_2), .IN3(na863_2), .IN4(~na864_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y110     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1491_4 ( .OUT(na1491_2), .IN1(1'b0), .IN2(1'b0), .IN3(na866_2), .IN4(na2749_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y94     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1492_1 ( .OUT(na1492_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2750_2), .IN6(1'b0), .IN7(1'b0), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x108y68     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1493_4 ( .OUT(na1493_2), .IN1(na875_2), .IN2(1'b0), .IN3(1'b0), .IN4(na2431_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y110     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1494_1 ( .OUT(na1494_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4216_2), .IN6(~na2752_1), .IN7(na863_2),
                      .IN8(na878_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y70     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1495_4 ( .OUT(na1495_2), .IN1(1'b0), .IN2(1'b0), .IN3(na881_1), .IN4(na2753_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x142y106     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1496_1 ( .OUT(na1496_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2434_2), .IN7(1'b0), .IN8(na884_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x138y100     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1497_4 ( .OUT(na1497_2), .IN1(na2435_2), .IN2(1'b0), .IN3(1'b0), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y107     80'h00_0060_00_0000_0C06_FF96
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1498_4 ( .OUT(na1498_2), .IN1(na2756_1), .IN2(na937_2), .IN3(~na938_1), .IN4(na936_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y110     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1499_1 ( .OUT(na1499_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2757_2), .IN6(~na943_2), .IN7(na938_1),
                      .IN8(na942_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y78     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1500_1 ( .OUT(na1500_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2758_1), .IN6(1'b0), .IN7(1'b0), .IN8(na948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x107y66     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1501_4 ( .OUT(na1501_2), .IN1(na2759_2), .IN2(1'b0), .IN3(na952_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y80     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1502_1 ( .OUT(na1502_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2440_2), .IN8(na955_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y88     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1503_1 ( .OUT(na1503_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na937_2), .IN7(~na2761_1), .IN8(na949_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y113     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1504_1 ( .OUT(na1504_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1480_1), .IN6(na2770_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x96y108     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1505_4 ( .OUT(na1505_2), .IN1(na2771_1), .IN2(na2739_1), .IN3(1'b0), .IN4(na263_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x94y77     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1506_1 ( .OUT(na1506_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2740_1), .IN7(na2772_2), .IN8(na275_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x87y116     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1507_4 ( .OUT(na1507_2), .IN1(na1483_2), .IN2(na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y73     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1508_1 ( .OUT(na1508_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1484_1), .IN6(1'b0), .IN7(1'b0), .IN8(na2774_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y79     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1509_4 ( .OUT(na1509_2), .IN1(na2775_1), .IN2(1'b0), .IN3(na298_1), .IN4(na2743_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x92y88     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1510_1 ( .OUT(na1510_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(1'b0), .IN7(na2776_1), .IN8(na2424_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x96y67     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1511_4 ( .OUT(na1511_2), .IN1(na312_1), .IN2(1'b0), .IN3(na2745_2), .IN4(na2777_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x119y116     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1512_4 ( .OUT(na1512_2), .IN1(na2778_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1488_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x137y107     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1513_1 ( .OUT(na1513_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na852_1), .IN6(na2779_1), .IN7(na2427_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y113     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1514_4 ( .OUT(na1514_2), .IN1(na2780_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1490_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y115     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1515_1 ( .OUT(na1515_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2781_1), .IN6(na4214_2), .IN7(na867_1),
                      .IN8(~na2749_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x133y98     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1516_4 ( .OUT(na1516_2), .IN1(na2750_2), .IN2(~na2782_2), .IN3(na873_1), .IN4(na864_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x106y67     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1517_4 ( .OUT(na1517_2), .IN1(na875_2), .IN2(1'b0), .IN3(na2783_1), .IN4(na2431_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x115y105     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1518_4 ( .OUT(na1518_2), .IN1(1'b0), .IN2(na2784_2), .IN3(1'b0), .IN4(na1494_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y78     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1519_1 ( .OUT(na1519_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2785_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1495_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y108     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1520_1 ( .OUT(na1520_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2786_2), .IN6(na2434_2), .IN7(1'b0), .IN8(na884_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x141y105     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1521_4 ( .OUT(na1521_2), .IN1(na2435_2), .IN2(na2787_1), .IN3(1'b0), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y116     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1522_1 ( .OUT(na1522_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2788_2), .IN6(1'b0), .IN7(na1498_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y110     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1523_1 ( .OUT(na1523_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1499_1), .IN7(na2789_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x118y87     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1524_4 ( .OUT(na1524_2), .IN1(~na2758_1), .IN2(~na2790_2), .IN3(na938_1), .IN4(na949_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x109y66     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1525_1 ( .OUT(na1525_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2759_2), .IN6(~na2791_1), .IN7(na953_1),
                      .IN8(na949_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y78     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1526_1 ( .OUT(na1526_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2792_2), .IN6(1'b0), .IN7(na2440_2), .IN8(na955_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y89     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1527_1 ( .OUT(na1527_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1503_1), .IN7(1'b0), .IN8(na2793_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x91y114     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1528_4 ( .OUT(na1528_2), .IN1(na1469_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2794_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x135y112     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1529_4 ( .OUT(na1529_2), .IN1(na4251_2), .IN2(~na2763_1), .IN3(~na3203_1), .IN4(na2795_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x108y115     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1530_4 ( .OUT(na1530_2), .IN1(1'b0), .IN2(na2796_2), .IN3(na1471_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x90y114     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1531_4 ( .OUT(na1531_2), .IN1(1'b0), .IN2(na1473_1), .IN3(1'b0), .IN4(na2797_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x97y116     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1532_4 ( .OUT(na1532_2), .IN1(na2798_2), .IN2(1'b0), .IN3(na1475_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y101     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1533_1 ( .OUT(na1533_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2799_1), .IN6(na1476_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x89y106     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1534_1 ( .OUT(na1534_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3208_2), .IN6(~na2768_2), .IN7(na2800_2),
                      .IN8(na1032_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y102     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1535_1 ( .OUT(na1535_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1478_1), .IN6(1'b0), .IN7(na2801_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x88y111     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1536_4 ( .OUT(na1536_2), .IN1(na1480_1), .IN2(na2770_2), .IN3(1'b0), .IN4(na2802_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x96y112     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1537_1 ( .OUT(na1537_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2803_1), .IN7(1'b0), .IN8(na1505_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y71     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1538_4 ( .OUT(na1538_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1506_1), .IN4(na2804_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y115     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1539_1 ( .OUT(na1539_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1483_2), .IN6(na2773_1), .IN7(1'b0), .IN8(na2805_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x94y81     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1540_4 ( .OUT(na1540_2), .IN1(na1484_1), .IN2(1'b0), .IN3(na2806_2), .IN4(na2774_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y86     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1541_1 ( .OUT(na1541_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1509_2), .IN8(na2807_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y90     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1542_1 ( .OUT(na1542_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(na2808_2), .IN7(~na2776_1),
                      .IN8(~na2424_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x91y67     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1543_1 ( .OUT(na1543_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1511_2), .IN8(na2809_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x121y116     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1544_4 ( .OUT(na1544_2), .IN1(na2778_2), .IN2(na2810_2), .IN3(1'b0), .IN4(na1488_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y108     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1545_1 ( .OUT(na1545_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na852_1), .IN6(~na2779_1), .IN7(~na2427_2),
                      .IN8(na2811_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y106     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1546_4 ( .OUT(na1546_2), .IN1(na2780_2), .IN2(na2812_2), .IN3(1'b0), .IN4(na1490_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x110y116     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1547_1 ( .OUT(na1547_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1515_1), .IN6(1'b0), .IN7(na2813_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y98     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1548_1 ( .OUT(na1548_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1516_2), .IN7(1'b0), .IN8(na2814_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x104y74     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1549_1 ( .OUT(na1549_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na875_2), .IN6(na2815_1), .IN7(~na2783_1),
                      .IN8(~na2431_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y109     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1550_1 ( .OUT(na1550_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2784_2), .IN7(na2816_2), .IN8(na1494_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x90y76     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1551_4 ( .OUT(na1551_2), .IN1(na2785_1), .IN2(na2817_1), .IN3(1'b0), .IN4(na1495_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x137y108     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1552_1 ( .OUT(na1552_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2786_2), .IN6(~na2434_2), .IN7(na2818_2),
                      .IN8(na884_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x140y101     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1553_4 ( .OUT(na1553_2), .IN1(~na2435_2), .IN2(~na2787_1), .IN3(na4229_2), .IN4(na2819_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y116     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1554_1 ( .OUT(na1554_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2788_2), .IN6(na2820_2), .IN7(na1498_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y112     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1555_4 ( .OUT(na1555_2), .IN1(1'b0), .IN2(na1499_1), .IN3(na2789_1), .IN4(na2821_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x115y87     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1556_4 ( .OUT(na1556_2), .IN1(1'b0), .IN2(na2822_2), .IN3(na1524_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x104y66     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1557_1 ( .OUT(na1557_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1525_1), .IN7(na2823_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x120y73     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1558_4 ( .OUT(na1558_2), .IN1(~na2792_2), .IN2(na2824_2), .IN3(~na2440_2), .IN4(na955_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y88     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1559_1 ( .OUT(na1559_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2825_1), .IN6(na1503_1), .IN7(1'b0), .IN8(na2793_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x98y111     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1560_4 ( .OUT(na1560_2), .IN1(na1469_1), .IN2(1'b0), .IN3(na2826_2), .IN4(na2794_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y110     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1561_1 ( .OUT(na1561_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1529_2), .IN7(1'b0), .IN8(na2827_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y116     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1562_1 ( .OUT(na1562_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2796_2), .IN7(na1471_1), .IN8(na2828_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x99y117     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1563_4 ( .OUT(na1563_2), .IN1(1'b0), .IN2(na1473_1), .IN3(na2829_1), .IN4(na2797_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y115     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1564_1 ( .OUT(na1564_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2798_2), .IN6(1'b0), .IN7(na1475_2), .IN8(na2830_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x91y94     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1565_4 ( .OUT(na1565_2), .IN1(na2799_1), .IN2(na1476_1), .IN3(1'b0), .IN4(na2831_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x87y100     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1566_4 ( .OUT(na1566_2), .IN1(1'b0), .IN2(na1534_1), .IN3(1'b0), .IN4(na2832_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y102     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1567_1 ( .OUT(na1567_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1478_1), .IN6(1'b0), .IN7(na2801_1), .IN8(na2833_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x89y110     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1568_4 ( .OUT(na1568_2), .IN1(na1480_1), .IN2(~na2770_2), .IN3(na2418_2), .IN4(~na2802_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x102y109     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1569_4 ( .OUT(na1569_2), .IN1(1'b0), .IN2(na2803_1), .IN3(na2419_1), .IN4(na1505_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y81     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1570_1 ( .OUT(na1570_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2420_2), .IN6(1'b0), .IN7(na1506_1), .IN8(na2804_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x88y113     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1571_4 ( .OUT(na1571_2), .IN1(na2421_1), .IN2(~na2773_1), .IN3(na4280_2), .IN4(~na2805_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y79     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1572_1 ( .OUT(na1572_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1484_1), .IN6(na2422_2), .IN7(~na2806_2),
                      .IN8(~na2774_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x101y83     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1573_4 ( .OUT(na1573_2), .IN1(1'b0), .IN2(na2423_1), .IN3(na1509_2), .IN4(na2807_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y90     80'h00_0018_00_0000_0666_9036
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1574_1 ( .OUT(na1574_1), .IN1(na308_1), .IN2(na2808_2), .IN3(1'b0), .IN4(~na2424_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na2776_1),
                      .IN8(na2424_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x92y67     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1575_1 ( .OUT(na1575_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2425_2), .IN6(1'b0), .IN7(na1511_2), .IN8(na2809_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x116y115     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1576_4 ( .OUT(na1576_2), .IN1(~na2778_2), .IN2(~na2810_2), .IN3(na2426_1), .IN4(na1488_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y107     80'h00_0018_00_0000_0666_A39A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1577_1 ( .OUT(na1577_1), .IN1(na852_1), .IN2(1'b0), .IN3(~na2427_2), .IN4(na2811_1), .IN5(1'b0), .IN6(~na2779_1), .IN7(na2427_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y106     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1578_1 ( .OUT(na1578_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2780_2), .IN6(~na2812_2), .IN7(na4281_2),
                      .IN8(na2428_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x109y116     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1579_1 ( .OUT(na1579_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1515_1), .IN6(1'b0), .IN7(na2813_1), .IN8(na2429_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y95     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1580_1 ( .OUT(na1580_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1516_2), .IN7(na2430_2), .IN8(na2814_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y73     80'h00_0018_00_0000_0666_60C6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1581_1 ( .OUT(na1581_1), .IN1(na875_2), .IN2(na2815_1), .IN3(1'b0), .IN4(na2431_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2783_1),
                      .IN8(~na2431_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x105y99     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1582_1 ( .OUT(na1582_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2432_1), .IN6(~na2784_2), .IN7(~na2816_2),
                      .IN8(na1494_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x91y69     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1583_4 ( .OUT(na1583_2), .IN1(~na2785_1), .IN2(~na2817_1), .IN3(na2433_2), .IN4(na1495_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y107     80'h00_0018_00_0000_0666_0963
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1584_1 ( .OUT(na1584_1), .IN1(1'b0), .IN2(~na2434_2), .IN3(na2818_2), .IN4(na884_1), .IN5(~na2786_2), .IN6(na2434_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y102     80'h00_0018_00_0000_0666_C9C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1585_1 ( .OUT(na1585_1), .IN1(~na2435_2), .IN2(1'b0), .IN3(1'b0), .IN4(na926_1), .IN5(na2435_1), .IN6(~na2787_1), .IN7(1'b0),
                      .IN8(na2819_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y114     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1586_1 ( .OUT(na1586_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2788_2), .IN6(~na2820_2), .IN7(na1498_2),
                      .IN8(na2436_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y110     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1587_4 ( .OUT(na1587_2), .IN1(na2437_1), .IN2(na1499_1), .IN3(~na2789_1), .IN4(~na2821_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x114y88     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1588_4 ( .OUT(na1588_2), .IN1(1'b0), .IN2(na2822_2), .IN3(na1524_2), .IN4(na2438_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x105y66     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1589_1 ( .OUT(na1589_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2439_2), .IN6(na1525_1), .IN7(na2823_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y80     80'h00_0018_00_0000_0666_A59C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1590_1 ( .OUT(na1590_1), .IN1(1'b0), .IN2(na2824_2), .IN3(~na2440_2), .IN4(na955_1), .IN5(~na2792_2), .IN6(1'b0), .IN7(na2440_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x90y77     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1591_4 ( .OUT(na1591_2), .IN1(~na2825_1), .IN2(na1503_1), .IN3(na2441_1), .IN4(~na2793_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x96y113     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1592_1 ( .OUT(na1592_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1469_1), .IN6(na2442_2), .IN7(~na2826_2),
                      .IN8(~na2794_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x133y108     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1593_4 ( .OUT(na1593_2), .IN1(na2443_1), .IN2(na1529_2), .IN3(1'b0), .IN4(na2827_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x113y115     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1594_1 ( .OUT(na1594_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2444_2), .IN6(~na2796_2), .IN7(na1471_1),
                      .IN8(~na2828_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x102y115     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1595_4 ( .OUT(na1595_2), .IN1(na2445_1), .IN2(na1473_1), .IN3(~na2829_1), .IN4(~na2797_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y111     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1596_1 ( .OUT(na1596_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2798_2), .IN6(na2446_2), .IN7(na1475_2),
                      .IN8(~na2830_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x87y96     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1597_4 ( .OUT(na1597_2), .IN1(~na2799_1), .IN2(na1476_1), .IN3(na4319_2), .IN4(~na2831_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y102     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1598_1 ( .OUT(na1598_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1534_1), .IN7(na2448_2), .IN8(na2832_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y99     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_1 ( .OUT(na1599_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1478_1), .IN6(~na4341_2), .IN7(na2449_1),
                      .IN8(~na2833_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y109     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1600_1 ( .OUT(na1600_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2834_2), .IN8(na4173_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x116y111     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1601_4 ( .OUT(na1601_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2835_2), .IN4(na263_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x98y78     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1602_1 ( .OUT(na1602_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2836_2), .IN6(1'b0), .IN7(1'b0), .IN8(na275_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x90y116     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1603_4 ( .OUT(na1603_2), .IN1(na2837_1), .IN2(1'b0), .IN3(na281_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x86y79     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1604_4 ( .OUT(na1604_2), .IN1(1'b0), .IN2(1'b0), .IN3(na293_1), .IN4(na2838_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x102y74     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1605_4 ( .OUT(na1605_2), .IN1(1'b0), .IN2(1'b0), .IN3(na298_1), .IN4(na2839_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x96y92     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1606_1 ( .OUT(na1606_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(na2464_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x100y66     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1607_4 ( .OUT(na1607_2), .IN1(na312_1), .IN2(na2841_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y112     80'h00_0060_00_0000_0C06_FF9A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1608_4 ( .OUT(na1608_2), .IN1(na808_2), .IN2(1'b0), .IN3(na848_1), .IN4(~na2842_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x142y106     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1609_4 ( .OUT(na1609_2), .IN1(na852_1), .IN2(na2467_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y110     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1610_1 ( .OUT(na1610_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na808_2), .IN6(~na2844_2), .IN7(na863_2), .IN8(~na864_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x124y105     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1611_4 ( .OUT(na1611_2), .IN1(na2845_1), .IN2(1'b0), .IN3(na866_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y89     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1612_1 ( .OUT(na1612_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2846_2), .IN6(1'b0), .IN7(1'b0), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x110y67     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1613_1 ( .OUT(na1613_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na875_2), .IN6(na2471_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x117y110     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1614_4 ( .OUT(na1614_2), .IN1(~na2848_1), .IN2(~na879_2), .IN3(na863_2), .IN4(na878_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x98y66     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1615_4 ( .OUT(na1615_2), .IN1(1'b0), .IN2(1'b0), .IN3(na881_1), .IN4(na2849_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y106     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1616_1 ( .OUT(na1616_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2474_2), .IN6(1'b0), .IN7(1'b0), .IN8(na884_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x141y104     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1617_4 ( .OUT(na1617_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2475_2), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y108     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1618_1 ( .OUT(na1618_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2852_1), .IN6(na937_2), .IN7(~na938_1), .IN8(na936_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x133y107     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1619_1 ( .OUT(na1619_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2853_2), .IN6(~na943_2), .IN7(na938_1),
                      .IN8(na942_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y78     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1620_1 ( .OUT(na1620_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2854_1), .IN7(1'b0), .IN8(na948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x107y67     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1621_4 ( .OUT(na1621_2), .IN1(1'b0), .IN2(na2855_2), .IN3(na952_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y82     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1622_4 ( .OUT(na1622_2), .IN1(na2480_2), .IN2(1'b0), .IN3(1'b0), .IN4(na955_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x102y84     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1623_1 ( .OUT(na1623_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na937_2), .IN7(na4231_2), .IN8(~na2857_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x96y116     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1624_1 ( .OUT(na1624_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na959_1), .IN6(na2858_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x136y110     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1625_4 ( .OUT(na1625_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2451_2), .IN4(na1003_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x111y116     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1626_1 ( .OUT(na1626_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2860_1), .IN6(na1014_2), .IN7(~na1016_1),
                      .IN8(na1013_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x113y115     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1627_4 ( .OUT(na1627_2), .IN1(~na4246_2), .IN2(na1020_1), .IN3(na1016_1), .IN4(na2861_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x99y113     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1628_4 ( .OUT(na1628_2), .IN1(na2862_1), .IN2(1'b0), .IN3(na1016_1), .IN4(na4254_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x100y80     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1629_4 ( .OUT(na1629_2), .IN1(na2863_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1029_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x99y94     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1630_1 ( .OUT(na1630_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2456_2), .IN7(1'b0), .IN8(na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y101     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1631_4 ( .OUT(na1631_2), .IN1(~na2865_1), .IN2(na1035_1), .IN3(na1030_1), .IN4(~na1015_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y114     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1632_1 ( .OUT(na1632_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1600_1), .IN8(na2279_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y112     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1633_1 ( .OUT(na1633_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2280_2), .IN7(na2835_2), .IN8(na263_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x94y74     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1634_4 ( .OUT(na1634_2), .IN1(na2836_2), .IN2(1'b0), .IN3(na4190_2), .IN4(na2281_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x87y113     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1635_4 ( .OUT(na1635_2), .IN1(na2282_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1603_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y91     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1636_1 ( .OUT(na1636_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2283_2), .IN6(1'b0), .IN7(na1604_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y80     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1637_1 ( .OUT(na1637_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2284_2), .IN7(na298_1), .IN8(na2839_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x90y88     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1638_4 ( .OUT(na1638_2), .IN1(na308_1), .IN2(na2464_2), .IN3(1'b0), .IN4(na2285_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x96y65     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1639_1 ( .OUT(na1639_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na312_1), .IN6(na2841_2), .IN7(na2286_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x109y113     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1640_4 ( .OUT(na1640_2), .IN1(1'b0), .IN2(na1608_2), .IN3(na2287_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x127y96     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1641_4 ( .OUT(na1641_2), .IN1(na852_1), .IN2(na2467_2), .IN3(1'b0), .IN4(na2288_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x130y108     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1642_1 ( .OUT(na1642_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2289_1), .IN7(1'b0), .IN8(na1610_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y111     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1643_1 ( .OUT(na1643_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2845_1), .IN6(~na2290_2), .IN7(na867_1),
                      .IN8(na864_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y100     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1644_1 ( .OUT(na1644_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2291_1), .IN6(na4342_2), .IN7(na873_1),
                      .IN8(na864_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x110y68     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1645_1 ( .OUT(na1645_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na875_2), .IN6(na2471_2), .IN7(na2292_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x104y108     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1646_1 ( .OUT(na1646_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1614_2), .IN7(1'b0), .IN8(na2293_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x94y66     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1647_4 ( .OUT(na1647_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2294_2), .IN4(na1615_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x134y108     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1648_4 ( .OUT(na1648_2), .IN1(na2474_2), .IN2(1'b0), .IN3(na2295_1), .IN4(na884_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y101     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1649_4 ( .OUT(na1649_2), .IN1(1'b0), .IN2(na2296_2), .IN3(na2475_2), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y114     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1650_1 ( .OUT(na1650_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2297_1), .IN7(1'b0), .IN8(na1618_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y106     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1651_4 ( .OUT(na1651_2), .IN1(na1619_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2298_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x113y90     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1652_1 ( .OUT(na1652_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2299_1), .IN6(~na2854_1), .IN7(na938_1),
                      .IN8(na949_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x104y66     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1653_4 ( .OUT(na1653_2), .IN1(~na2300_2), .IN2(na2855_2), .IN3(na953_1), .IN4(na949_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y81     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1654_4 ( .OUT(na1654_2), .IN1(na2480_2), .IN2(na2301_1), .IN3(1'b0), .IN4(na955_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x94y76     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1655_4 ( .OUT(na1655_2), .IN1(1'b0), .IN2(na2302_2), .IN3(1'b0), .IN4(na1623_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x92y116     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1656_1 ( .OUT(na1656_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2303_1), .IN8(na1624_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y111     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1657_1 ( .OUT(na1657_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2304_2), .IN7(na2451_2), .IN8(na1003_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x105y115     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1658_4 ( .OUT(na1658_2), .IN1(na2305_1), .IN2(na1626_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x104y115     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1659_4 ( .OUT(na1659_2), .IN1(na1627_2), .IN2(na2306_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y111     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1660_1 ( .OUT(na1660_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1628_2), .IN6(na2307_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x93y95     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1661_4 ( .OUT(na1661_2), .IN1(na2863_2), .IN2(~na2308_2), .IN3(na1030_1), .IN4(na4253_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x106y95     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1662_4 ( .OUT(na1662_2), .IN1(na2309_1), .IN2(na2456_2), .IN3(1'b0), .IN4(na1032_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x87y93     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1663_4 ( .OUT(na1663_2), .IN1(na2310_2), .IN2(1'b0), .IN3(na1631_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y111     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1664_1 ( .OUT(na1664_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2866_2), .IN7(na1600_1), .IN8(na2279_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x104y114     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1665_4 ( .OUT(na1665_2), .IN1(na2867_1), .IN2(na1633_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y79     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1666_1 ( .OUT(na1666_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2868_2), .IN8(na1634_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x88y116     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1667_4 ( .OUT(na1667_2), .IN1(na2282_2), .IN2(na2869_1), .IN3(1'b0), .IN4(na1603_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y89     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1668_1 ( .OUT(na1668_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2283_2), .IN6(na2870_2), .IN7(na1604_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y72     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1669_4 ( .OUT(na1669_2), .IN1(1'b0), .IN2(na1637_1), .IN3(na2871_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y88     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1670_4 ( .OUT(na1670_2), .IN1(na308_1), .IN2(~na2464_2), .IN3(na2872_1), .IN4(~na2285_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x95y66     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1671_4 ( .OUT(na1671_2), .IN1(1'b0), .IN2(na2873_1), .IN3(na1639_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x114y115     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1672_4 ( .OUT(na1672_2), .IN1(na2874_2), .IN2(na1608_2), .IN3(na2287_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x140y106     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1673_4 ( .OUT(na1673_2), .IN1(na852_1), .IN2(~na2467_2), .IN3(na2875_1), .IN4(~na2288_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y108     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1674_1 ( .OUT(na1674_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2289_1), .IN7(na2876_2), .IN8(na1610_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x117y116     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1675_4 ( .OUT(na1675_2), .IN1(na1643_1), .IN2(1'b0), .IN3(na2877_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y102     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1676_4 ( .OUT(na1676_2), .IN1(1'b0), .IN2(na1644_1), .IN3(na2878_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x105y67     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1677_4 ( .OUT(na1677_2), .IN1(na2879_1), .IN2(~na2471_2), .IN3(~na2292_2), .IN4(na4215_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x105y103     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1678_4 ( .OUT(na1678_2), .IN1(na2880_2), .IN2(na1614_2), .IN3(1'b0), .IN4(na2293_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x92y66     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1679_1 ( .OUT(na1679_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2881_1), .IN7(na2294_2), .IN8(na1615_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y108     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1680_1 ( .OUT(na1680_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2474_2), .IN6(na2882_2), .IN7(~na2295_1),
                      .IN8(na884_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y103     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1681_4 ( .OUT(na1681_2), .IN1(na2883_1), .IN2(~na2296_2), .IN3(~na2475_2), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x119y113     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1682_4 ( .OUT(na1682_2), .IN1(na2884_2), .IN2(na2297_1), .IN3(1'b0), .IN4(na1618_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x133y109     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1683_1 ( .OUT(na1683_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1619_1), .IN6(na2885_1), .IN7(1'b0), .IN8(na2298_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x106y85     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1684_1 ( .OUT(na1684_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1652_1), .IN7(na2886_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x102y65     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1685_1 ( .OUT(na1685_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2887_1), .IN8(na1653_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y81     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1686_1 ( .OUT(na1686_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2480_2), .IN6(~na2301_1), .IN7(na2888_2),
                      .IN8(na955_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x90y80     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1687_4 ( .OUT(na1687_2), .IN1(1'b0), .IN2(na2302_2), .IN3(na2889_1), .IN4(na1623_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x94y116     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1688_1 ( .OUT(na1688_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2890_2), .IN7(na2303_1), .IN8(na1624_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x135y109     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1689_4 ( .OUT(na1689_2), .IN1(na2891_1), .IN2(~na2304_2), .IN3(~na2451_2), .IN4(na1003_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x106y116     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1690_4 ( .OUT(na1690_2), .IN1(na2305_1), .IN2(na1626_1), .IN3(na2892_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x103y115     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1691_1 ( .OUT(na1691_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1627_2), .IN6(na2306_2), .IN7(na2893_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y110     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1692_1 ( .OUT(na1692_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1628_2), .IN6(na2307_1), .IN7(na2894_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x87y89     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1693_4 ( .OUT(na1693_2), .IN1(na1661_2), .IN2(1'b0), .IN3(na2895_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x102y107     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1694_4 ( .OUT(na1694_2), .IN1(~na2309_1), .IN2(~na2456_2), .IN3(na2896_2), .IN4(na1032_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y95     80'h00_0018_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1695_1 ( .OUT(na1695_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2310_2), .IN6(na2897_1), .IN7(na1631_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y110     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1696_1 ( .OUT(na1696_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2458_2), .IN6(~na2866_2), .IN7(na1600_1),
                      .IN8(~na2279_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x113y114     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1697_4 ( .OUT(na1697_2), .IN1(na2459_1), .IN2(na1633_1), .IN3(na4343_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x104y82     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1698_1 ( .OUT(na1698_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4326_2), .IN6(1'b0), .IN7(na2868_2), .IN8(na1634_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x91y115     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1699_4 ( .OUT(na1699_2), .IN1(~na2282_2), .IN2(~na2869_1), .IN3(na2461_1), .IN4(na1603_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y90     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1700_1 ( .OUT(na1700_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2462_2), .IN6(~na2870_2), .IN7(na1604_2),
                      .IN8(~na4305_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x88y75     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1701_4 ( .OUT(na1701_2), .IN1(na2463_1), .IN2(na1637_1), .IN3(na2871_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y93     80'h00_0018_00_0000_0666_39AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1702_1 ( .OUT(na1702_1), .IN1(1'b0), .IN2(na2464_1), .IN3(na2872_1), .IN4(1'b0), .IN5(na308_1), .IN6(~na2464_2), .IN7(1'b0),
                      .IN8(~na2285_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x94y66     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1703_1 ( .OUT(na1703_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2873_1), .IN7(na1639_1), .IN8(na4328_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x115y116     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1704_1 ( .OUT(na1704_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2874_2), .IN6(na1608_2), .IN7(~na2287_1),
                      .IN8(na2466_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x141y107     80'h00_0018_00_0000_0666_39AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1705_1 ( .OUT(na1705_1), .IN1(1'b0), .IN2(na2467_1), .IN3(na2875_1), .IN4(1'b0), .IN5(na852_1), .IN6(~na2467_2), .IN7(1'b0),
                      .IN8(~na2288_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x132y107     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1706_4 ( .OUT(na1706_2), .IN1(na2468_2), .IN2(~na2289_1), .IN3(~na2876_2), .IN4(na1610_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x115y114     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1707_4 ( .OUT(na1707_2), .IN1(na1643_1), .IN2(na2469_1), .IN3(na2877_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y99     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1708_1 ( .OUT(na1708_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1644_1), .IN7(na2878_2), .IN8(na2470_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y68     80'h00_0018_00_0000_0666_5906
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1709_1 ( .OUT(na1709_1), .IN1(na875_2), .IN2(na2471_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2879_1), .IN6(~na2471_2), .IN7(~na2292_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x112y100     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1710_4 ( .OUT(na1710_2), .IN1(~na2880_2), .IN2(na1614_2), .IN3(na2472_1), .IN4(~na2293_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x95y67     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1711_1 ( .OUT(na1711_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2473_1), .IN6(~na2881_1), .IN7(~na2294_2),
                      .IN8(na1615_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x133y110     80'h00_0018_00_0000_0666_9506
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1712_1 ( .OUT(na1712_1), .IN1(na2474_1), .IN2(na2882_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2474_2), .IN6(1'b0), .IN7(~na2295_1),
                      .IN8(na884_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x137y97     80'h00_0018_00_0000_0666_635A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1713_1 ( .OUT(na1713_1), .IN1(na2883_1), .IN2(1'b0), .IN3(~na2475_2), .IN4(1'b0), .IN5(1'b0), .IN6(~na2296_2), .IN7(na2475_1),
                      .IN8(na926_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x118y114     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1714_4 ( .OUT(na1714_2), .IN1(~na2884_2), .IN2(~na2297_1), .IN3(na2476_1), .IN4(na1618_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y99     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1715_1 ( .OUT(na1715_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1619_1), .IN6(~na2885_1), .IN7(na2477_2),
                      .IN8(~na2298_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x109y87     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1716_4 ( .OUT(na1716_2), .IN1(na2478_1), .IN2(na1652_1), .IN3(na2886_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x102y67     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1717_1 ( .OUT(na1717_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2479_2), .IN7(na2887_1), .IN8(na1653_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y84     80'h00_0018_00_0000_0666_6905
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1718_1 ( .OUT(na1718_1), .IN1(~na2480_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2480_1), .IN6(~na2301_1), .IN7(na2888_2),
                      .IN8(na955_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y83     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1719_1 ( .OUT(na1719_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2481_1), .IN6(~na2302_2), .IN7(~na2889_1),
                      .IN8(na1623_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x94y115     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1720_4 ( .OUT(na1720_2), .IN1(na2450_2), .IN2(~na2890_2), .IN3(~na2303_1), .IN4(na1624_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y106     80'h00_0018_00_0000_0666_93AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1721_1 ( .OUT(na1721_1), .IN1(na2891_1), .IN2(1'b0), .IN3(na2451_1), .IN4(1'b0), .IN5(1'b0), .IN6(~na2304_2), .IN7(~na2451_2),
                      .IN8(na1003_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x108y116     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1722_1 ( .OUT(na1722_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2305_1), .IN6(na1626_1), .IN7(na2452_1),
                      .IN8(~na4344_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x104y116     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1723_1 ( .OUT(na1723_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1627_2), .IN6(~na2306_2), .IN7(~na2893_1),
                      .IN8(na2453_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y110     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1724_4 ( .OUT(na1724_2), .IN1(na1628_2), .IN2(~na2307_1), .IN3(~na2894_2), .IN4(na2454_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y91     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1725_4 ( .OUT(na1725_2), .IN1(na1661_2), .IN2(1'b0), .IN3(na2455_2), .IN4(na4345_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x93y103     80'h00_0018_00_0000_0666_C6AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1726_1 ( .OUT(na1726_1), .IN1(1'b0), .IN2(na2456_1), .IN3(na2896_2), .IN4(1'b0), .IN5(~na2309_1), .IN6(~na2456_2), .IN7(1'b0),
                      .IN8(na1032_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x91y95     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1727_1 ( .OUT(na1727_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2310_2), .IN6(~na2897_1), .IN7(na1631_2),
                      .IN8(na4325_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x109y71     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1728_1 ( .OUT(na1728_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4347_2), .IN6(na1729_1), .IN7(na2953_1),
                      .IN8(~na2969_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x113y70     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1729_1 ( .OUT(na1729_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2957_2), .IN6(1'b0), .IN7(na2970_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x113y69     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1730_1 ( .OUT(na1730_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2955_1), .IN6(na1729_1), .IN7(na1731_1),
                      .IN8(~na1732_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y69     80'h00_0018_00_0000_0C66_5C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1731_1 ( .OUT(na1731_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2946_1), .IN7(~na2953_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x118y70     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1732_4 ( .OUT(na1732_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2963_2), .IN4(na2971_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y70     80'h00_0018_00_0000_0666_6C06
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1733_1 ( .OUT(na1733_1), .IN1(na4348_2), .IN2(na2965_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2956_1), .IN7(na2964_1),
                      .IN8(na2971_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y71     80'h00_0018_00_0000_0666_5669
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1735_1 ( .OUT(na1735_1), .IN1(na2957_1), .IN2(~na2965_2), .IN3(~na2953_1), .IN4(~na4349_2), .IN5(na2957_2), .IN6(na2965_1),
                      .IN7(~na2953_2), .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y68     80'h00_0018_00_0000_0666_9C96
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1737_1 ( .OUT(na1737_1), .IN1(na2957_2), .IN2(na2966_1), .IN3(na2953_1), .IN4(~na2949_1), .IN5(1'b0), .IN6(na2966_2), .IN7(na2953_2),
                      .IN8(~na2949_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y66     80'h00_0018_00_0000_0666_AA59
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1739_1 ( .OUT(na1739_1), .IN1(na2959_1), .IN2(~na2966_2), .IN3(~na2950_2), .IN4(1'b0), .IN5(na2959_2), .IN6(1'b0), .IN7(na2967_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y65     80'h00_0018_00_0000_0666_633A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1741_1 ( .OUT(na1741_1), .IN1(na2959_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na2968_2), .IN5(1'b0), .IN6(~na2976_1), .IN7(na2967_2),
                      .IN8(na2968_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y66     80'h00_0018_00_0000_0666_C909
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1743_1 ( .OUT(na1743_1), .IN1(~na2961_1), .IN2(na2976_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2957_2), .IN6(na2976_2), .IN7(1'b0),
                      .IN8(na2969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x113y69     80'h00_0060_00_0000_0C06_FF96
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1745_4 ( .OUT(na1745_2), .IN1(na2961_1), .IN2(na4352_2), .IN3(na1731_1), .IN4(~na2969_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x116y69     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1746_1 ( .OUT(na1746_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1747_1), .IN6(~na2956_2), .IN7(na1731_1),
                      .IN8(na1732_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x115y69     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1747_1 ( .OUT(na1747_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2961_1), .IN6(na2946_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y69     80'h00_0018_00_0000_0666_09A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1748_1 ( .OUT(na1748_1), .IN1(na2955_1), .IN2(~na2965_2), .IN3(na2964_1), .IN4(1'b0), .IN5(na2961_2), .IN6(~na2956_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x111y70     80'h00_0018_00_0000_0666_69A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1750_1 ( .OUT(na1750_1), .IN1(~na2961_2), .IN2(na2965_1), .IN3(na2953_2), .IN4(1'b0), .IN5(na2961_1), .IN6(~na2956_1), .IN7(na2953_1),
                      .IN8(na2949_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y67     80'h00_0018_00_0000_0666_A699
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1752_1 ( .OUT(na1752_1), .IN1(na2961_1), .IN2(~na2966_2), .IN3(na2950_2), .IN4(~na2949_1), .IN5(na2957_1), .IN6(na2966_1),
                      .IN7(na2953_1), .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x115y66     80'h00_0018_00_0000_0666_6059
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1754_1 ( .OUT(na1754_1), .IN1(~na2959_2), .IN2(na4350_2), .IN3(~na2967_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2950_2),
                      .IN8(na2949_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y67     80'h00_0018_00_0000_0666_660C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1756_1 ( .OUT(na1756_1), .IN1(1'b0), .IN2(na2976_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2959_1), .IN6(na2976_1), .IN7(na2967_2),
                      .IN8(na2968_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x113y68     80'h00_0018_00_0000_0666_65C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1758_1 ( .OUT(na1758_1), .IN1(1'b0), .IN2(~na2976_2), .IN3(1'b0), .IN4(na2969_1), .IN5(~na2957_2), .IN6(1'b0), .IN7(na2953_1),
                      .IN8(na2968_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x116y69     80'h00_0060_00_0000_0C06_FF96
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1760_4 ( .OUT(na1760_2), .IN1(na1747_1), .IN2(na2946_1), .IN3(~na2970_2), .IN4(na2969_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y70     80'h00_0018_00_0000_0666_C9C6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1761_1 ( .OUT(na1761_1), .IN1(na1747_1), .IN2(na2956_2), .IN3(1'b0), .IN4(na2969_2), .IN5(~na2955_1), .IN6(na4351_2), .IN7(1'b0),
                      .IN8(na2971_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y69     80'h00_0018_00_0000_0666_A606
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1763_1 ( .OUT(na1763_1), .IN1(~na2955_1), .IN2(~na2965_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2961_2), .IN6(na2956_1), .IN7(na2963_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y70     80'h00_0018_00_0000_0666_6965
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1765_1 ( .OUT(na1765_1), .IN1(~na2957_1), .IN2(1'b0), .IN3(na2953_2), .IN4(na2969_1), .IN5(na2961_1), .IN6(~na2956_1), .IN7(na2964_1),
                      .IN8(na2949_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y68     80'h00_0018_00_0000_0666_C699
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1767_1 ( .OUT(na1767_1), .IN1(na2961_1), .IN2(~na2965_1), .IN3(na2950_2), .IN4(~na2949_2), .IN5(na2957_1), .IN6(na2966_2),
                      .IN7(1'b0), .IN8(na2969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y65     80'h00_0018_00_0000_0666_563A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1769_1 ( .OUT(na1769_1), .IN1(na2959_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na2949_2), .IN5(na2959_2), .IN6(na2966_1), .IN7(~na2967_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y66     80'h00_0018_00_0000_0666_9C09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1770_1 ( .OUT(na1770_1), .IN1(~na2959_1), .IN2(na2976_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2976_1), .IN7(na2967_1),
                      .IN8(~na2968_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y67     80'h00_0018_00_0000_0666_CA6A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1771_1 ( .OUT(na1771_1), .IN1(na2957_2), .IN2(1'b0), .IN3(~na2953_1), .IN4(~na2968_2), .IN5(na2961_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na2968_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y72     80'h00_0018_00_0000_0666_36C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1773_1 ( .OUT(na1773_1), .IN1(1'b0), .IN2(~na2946_2), .IN3(1'b0), .IN4(na2969_1), .IN5(na2957_2), .IN6(na2946_1), .IN7(1'b0),
                      .IN8(~na2969_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y70     80'h00_0018_00_0000_0666_C69C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1775_1 ( .OUT(na1775_1), .IN1(1'b0), .IN2(na2956_2), .IN3(~na2963_2), .IN4(na2969_2), .IN5(na2955_1), .IN6(na1729_1), .IN7(1'b0),
                      .IN8(na2969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x119y71     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1776_4 ( .OUT(na1776_2), .IN1(~na2961_2), .IN2(~na2956_1), .IN3(na2964_1), .IN4(na1732_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y72     80'h00_0018_00_0000_0666_69C9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1777_1 ( .OUT(na1777_1), .IN1(~na2957_2), .IN2(na2965_2), .IN3(1'b0), .IN4(na2949_1), .IN5(~na2957_1), .IN6(na2965_1), .IN7(na2964_1),
                      .IN8(na2969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x111y69     80'h00_0018_00_0000_0666_6963
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1779_1 ( .OUT(na1779_1), .IN1(1'b0), .IN2(~na2965_1), .IN3(na2950_2), .IN4(na2969_1), .IN5(na2957_2), .IN6(~na2966_1), .IN7(na2953_2),
                      .IN8(na2949_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x115y68     80'h00_0018_00_0000_0666_565C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1781_1 ( .OUT(na1781_1), .IN1(1'b0), .IN2(na2966_1), .IN3(~na2967_2), .IN4(1'b0), .IN5(na2959_1), .IN6(na2966_2), .IN7(~na2967_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y67     80'h00_0018_00_0000_0666_3C9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1783_1 ( .OUT(na1783_1), .IN1(na2959_2), .IN2(1'b0), .IN3(na2967_1), .IN4(~na2968_1), .IN5(1'b0), .IN6(na2976_2), .IN7(1'b0),
                      .IN8(~na2968_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x111y68     80'h00_0018_00_0000_0666_63C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1784_1 ( .OUT(na1784_1), .IN1(~na2961_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2969_1), .IN5(1'b0), .IN6(~na2976_1), .IN7(na2953_1),
                      .IN8(na2968_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y118     80'h00_0018_00_0000_0666_C6AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1797_1 ( .OUT(na1797_1), .IN1(1'b0), .IN2(na225_1), .IN3(na222_2), .IN4(1'b0), .IN5(~na223_1), .IN6(~na224_1), .IN7(1'b0),
                      .IN8(na4103_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y115     80'h00_0018_00_0000_0666_ACC9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1799_1 ( .OUT(na1799_1), .IN1(na228_2), .IN2(~na4104_1), .IN3(1'b0), .IN4(na4105_2), .IN5(1'b0), .IN6(na229_1), .IN7(na4177_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y115     80'h00_0018_00_0040_0A79_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1800_1 ( .OUT(na1800_1), .IN1(~na223_1), .IN2(1'b1), .IN3(1'b1), .IN4(na227_1), .IN5(~na226_1), .IN6(na253_2), .IN7(na236_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y114     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1801_1 ( .OUT(na1801_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na237_1), .IN6(1'b0), .IN7(na1800_1), .IN8(na238_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y90     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1803_1 ( .OUT(na1803_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2898_2),
                      .IN8(~na2359_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x109y73     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1804_4 ( .OUT(na1804_2), .IN1(na4109_2), .IN2(na57_2), .IN3(~na260_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x108y86     80'h00_0018_00_0040_0C4A_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1805_1 ( .OUT(na1805_1), .IN1(1'b0), .IN2(na262_2), .IN3(1'b1), .IN4(na4110_1), .IN5(1'b1), .IN6(na57_2), .IN7(~na26_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x108y76     80'h00_0018_00_0040_0C5A_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1806_1 ( .OUT(na1806_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(na4111_2), .IN5(na1804_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1805_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y92     80'h00_0018_00_0040_0A3F_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1808_1 ( .OUT(na1808_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(~na2360_2), .IN6(~na2899_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x115y79     80'h00_0018_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1809_1 ( .OUT(na1809_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4114_1), .IN6(na57_2), .IN7(1'b0), .IN8(~na272_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x116y86     80'h00_0018_00_0040_0C25_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1810_1 ( .OUT(na1810_1), .IN1(na4115_1), .IN2(1'b1), .IN3(na274_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na57_2), .IN7(na26_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x112y80     80'h00_0018_00_0040_0C5A_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1811_1 ( .OUT(na1811_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(na4116_1), .IN5(na1809_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1810_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y85     80'h00_0018_00_0040_0A5F_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1813_1 ( .OUT(na1813_1), .IN1(1'b1), .IN2(na4164_2), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2900_2), .IN6(1'b1), .IN7(~na2361_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x111y67     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1814_4 ( .OUT(na1814_2), .IN1(na4119_1), .IN2(na57_2), .IN3(~na278_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x112y83     80'h00_0018_00_0040_0C1A_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1815_1 ( .OUT(na1815_1), .IN1(1'b1), .IN2(na4120_1), .IN3(1'b0), .IN4(na280_1), .IN5(1'b1), .IN6(na57_2), .IN7(na26_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x110y72     80'h00_0018_00_0040_0C5A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1816_1 ( .OUT(na1816_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(na4121_2), .IN5(na1814_2), .IN6(1'b1), .IN7(na1815_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y86     80'h00_0018_00_0040_0A3F_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1818_1 ( .OUT(na1818_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(~na2363_1), .IN6(~na2902_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x111y71     80'h00_0018_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1819_1 ( .OUT(na1819_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4124_2), .IN6(na57_2), .IN7(~na295_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x104y79     80'h00_0018_00_0040_0C1A_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1820_1 ( .OUT(na1820_1), .IN1(1'b1), .IN2(na4125_1), .IN3(1'b0), .IN4(na297_2), .IN5(1'b1), .IN6(na57_2), .IN7(na26_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y70     80'h00_0018_00_0040_0C5A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1821_1 ( .OUT(na1821_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(na4126_2), .IN5(na1819_1), .IN6(1'b1), .IN7(na1820_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y86     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1823_1 ( .OUT(na1823_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na19_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2365_1),
                      .IN8(~na2904_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x107y69     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1824_4 ( .OUT(na1824_2), .IN1(na4129_2), .IN2(na57_2), .IN3(~na309_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x108y78     80'h00_0018_00_0040_0C1A_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1825_1 ( .OUT(na1825_1), .IN1(1'b1), .IN2(na4130_1), .IN3(1'b0), .IN4(na311_1), .IN5(1'b1), .IN6(na57_2), .IN7(na26_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y72     80'h00_0018_00_0040_0C5A_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1826_1 ( .OUT(na1826_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(na4131_2), .IN5(na1824_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1825_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y82     80'h00_0018_00_0040_0A3F_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1828_1 ( .OUT(na1828_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(na19_1), .IN5(~na2905_1), .IN6(~na2366_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x109y66     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1829_4 ( .OUT(na1829_2), .IN1(na4134_2), .IN2(na57_2), .IN3(~na313_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x102y76     80'h00_0018_00_0040_0C1A_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1830_1 ( .OUT(na1830_1), .IN1(1'b1), .IN2(na4135_1), .IN3(1'b0), .IN4(na315_1), .IN5(1'b1), .IN6(na57_2), .IN7(na26_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x110y69     80'h00_0018_00_0040_0C5A_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1831_1 ( .OUT(na1831_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(na4136_1), .IN5(1'b1), .IN6(na1829_2), .IN7(1'b1), .IN8(na1830_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x149y113     80'h00_0018_00_0040_0AFA_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1832_1 ( .OUT(na1832_1), .IN1(na817_1), .IN2(1'b1), .IN3(~na4201_2), .IN4(1'b1), .IN5(na4200_2), .IN6(~na813_1), .IN7(na812_2),
                      .IN8(~na4199_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x150y115     80'h00_0060_00_0000_0C06_FFE5
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1833_4 ( .OUT(na1833_2), .IN1(na1832_1), .IN2(1'b1), .IN3(~na815_2), .IN4(~na3704_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x145y115     80'h00_0018_00_0000_0C66_AEFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1834_1 ( .OUT(na1834_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4203_2), .IN6(~na818_1), .IN7(~na1833_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x144y116     80'h00_0018_00_0040_0A7C_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1835_1 ( .OUT(na1835_1), .IN1(na823_1), .IN2(1'b1), .IN3(~na815_2), .IN4(1'b1), .IN5(na4359_2), .IN6(na813_1), .IN7(~na4401_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y114     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1836_4 ( .OUT(na1836_2), .IN1(1'b0), .IN2(na829_1), .IN3(na828_2), .IN4(na1835_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x150y100     80'h00_0018_00_0040_0C49_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1837_1 ( .OUT(na1837_1), .IN1(na4367_2), .IN2(1'b0), .IN3(1'b1), .IN4(na3031_2), .IN5(1'b1), .IN6(na4371_2), .IN7(~na3030_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y97     80'h00_0018_00_0040_0A72_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1838_1 ( .OUT(na1838_1), .IN1(1'b1), .IN2(na4371_2), .IN3(1'b1), .IN4(na3033_1), .IN5(na3027_1), .IN6(~na4368_2), .IN7(na4141_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x145y101     80'h00_0018_00_0000_0666_F537
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1839_1 ( .OUT(na1839_1), .IN1(na892_2), .IN2(na894_2), .IN3(1'b1), .IN4(na1837_1), .IN5(na1838_1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x147y103     80'h00_0018_00_0000_0C66_3D00
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1840_1 ( .OUT(na1840_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na892_2), .IN6(~na3748_2), .IN7(1'b1), .IN8(na3031_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x148y108     80'h00_0018_00_0000_0666_EABA
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1841_1 ( .OUT(na1841_1), .IN1(~na1840_1), .IN2(1'b1), .IN3(~na3026_2), .IN4(na893_2), .IN5(~na899_1), .IN6(1'b1), .IN7(~na897_1),
                      .IN8(~na891_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x149y111     80'h00_0018_00_0040_0AD2_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1842_1 ( .OUT(na1842_1), .IN1(1'b1), .IN2(na4221_2), .IN3(1'b1), .IN4(na893_2), .IN5(na4146_1), .IN6(1'b1), .IN7(na3026_2),
                      .IN8(na891_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y106     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1843_4 ( .OUT(na1843_2), .IN1(na1842_1), .IN2(na902_1), .IN3(na901_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y111     80'h00_0060_00_0000_0C06_FF3A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1844_4 ( .OUT(na1844_2), .IN1(na4147_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na968_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x139y117     80'h00_0018_00_0000_0C66_E500
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1845_1 ( .OUT(na1845_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1844_2), .IN6(1'b1), .IN7(~na966_2), .IN8(~na3781_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x140y115     80'h00_0060_00_0000_0C06_FFEA
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1846_4 ( .OUT(na1846_2), .IN1(~na1845_1), .IN2(1'b1), .IN3(~na4236_2), .IN4(~na969_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y118     80'h00_0018_00_0040_0A78_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1847_1 ( .OUT(na1847_1), .IN1(1'b1), .IN2(na974_1), .IN3(~na966_2), .IN4(1'b1), .IN5(na3034_2), .IN6(na964_1), .IN7(na4151_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y116     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1848_1 ( .OUT(na1848_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na980_1), .IN6(na1847_1), .IN7(1'b0), .IN8(na979_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y68     80'h00_0018_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1849_1 ( .OUT(na1849_1), .IN1(1'b1), .IN2(1'b1), .IN3(na3151_2), .IN4(1'b1), .IN5(1'b0), .IN6(na57_2), .IN7(1'b0), .IN8(na1948_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y66     80'h00_0018_00_0040_0AB4_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1850_1 ( .OUT(na1850_1), .IN1(~na4381_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3150_2), .IN5(na4153_1), .IN6(na4152_2), .IN7(1'b1),
                      .IN8(na4416_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y92     80'h00_0078_00_0020_0C66_3303
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1852_1 ( .OUT(na1852_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1941_2), .IN7(1'b1), .IN8(~na1946_2),
                      .CINX(1'b0), .CINY1(na1859_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1852_4 ( .OUT(na1852_2), .COUTY1(na1852_4), .IN1(1'b1), .IN2(~na1941_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1941_2),
                      .IN7(1'b1), .IN8(~na1946_2), .CINX(1'b0), .CINY1(na1859_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y93     80'h00_0078_00_0020_0C66_5050
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1854_1 ( .OUT(na1854_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1943_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1852_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1854_4 ( .OUT(na1854_2), .COUTY1(na1854_4), .IN1(1'b0), .IN2(1'b0), .IN3(~na1943_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(~na1943_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1852_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y94     80'h00_0078_00_0020_0C66_0505
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1856_1 ( .OUT(na1856_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1945_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1854_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1856_4 ( .OUT(na1856_2), .COUTY1(na1856_4), .IN1(~na1945_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1945_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1854_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x143y95     80'h00_0018_00_0010_0666_0030
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1858_1 ( .OUT(na1858_1), .COUTY1(na1858_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1946_1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1856_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x143y91     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1859_2 ( .OUT(na1859_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1859_6 ( .COUTY1(na1859_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1859_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x89y112     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1860_1 ( .OUT(na1860_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1935_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1934_2),
                      .CINX(1'b0), .CINY1(na1865_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1860_4 ( .OUT(na1860_2), .COUTY1(na1860_4), .IN1(na1935_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1935_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na1934_2), .CINX(1'b0), .CINY1(na1865_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y113     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1862_1 ( .OUT(na1862_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1937_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1860_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1862_4 ( .OUT(na1862_2), .COUTY1(na1862_4), .IN1(1'b1), .IN2(na1937_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1937_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1860_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x89y114     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1864_1 ( .OUT(na1864_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1938_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1862_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x89y111     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1865_2 ( .OUT(na1865_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1865_6 ( .COUTY1(na1865_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1865_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x145y85     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1866_1 ( .OUT(na1866_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1929_1), .IN7(na1930_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1870_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1866_4 ( .OUT(na1866_2), .COUTY1(na1866_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1930_1), .IN4(1'b1), .IN5(1'b1), .IN6(na1929_1),
                      .IN7(na1930_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1870_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x145y86     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1868_1 ( .OUT(na1868_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1932_2),
                      .CINX(1'b0), .CINY1(na1866_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1868_4 ( .OUT(na1868_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1932_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1932_2),
                      .CINX(1'b0), .CINY1(na1866_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x145y84     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1870_2 ( .OUT(na1870_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1870_6 ( .COUTY1(na1870_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1870_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x124y74     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1871_1 ( .OUT(na1871_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2416_2), .IN7(na4309_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1874_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1871_4 ( .OUT(na1871_2), .COUTY1(na1871_4), .IN1(1'b1), .IN2(na2416_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2416_2),
                      .IN7(na4309_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1874_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x124y75     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1873_1 ( .OUT(na1873_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2417_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1871_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x124y73     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1874_2 ( .OUT(na1874_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1874_6 ( .COUTY1(na1874_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1874_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x89y72     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1876_1 ( .OUT(na1876_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4386_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3173_1),
                      .CINX(1'b0), .CINY1(na1885_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1876_4 ( .OUT(na1876_2), .COUTY1(na1876_4), .IN1(na3175_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4386_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na3173_1), .CINX(1'b0), .CINY1(na1885_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y73     80'h00_0078_00_0020_0C66_0C0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1878_1 ( .OUT(na1878_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3176_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1876_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1878_4 ( .OUT(na1878_2), .COUTY1(na1878_4), .IN1(na3175_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3176_1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1876_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y74     80'h00_0078_00_0020_0C66_0AC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1880_1 ( .OUT(na1880_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3178_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1878_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1880_4 ( .OUT(na1880_2), .COUTY1(na1880_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3182_2), .IN5(na3178_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1878_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y75     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1882_1 ( .OUT(na1882_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3180_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1880_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1882_4 ( .OUT(na1882_2), .COUTY1(na1882_4), .IN1(1'b1), .IN2(na3181_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3180_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1880_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y76     80'h00_0078_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1884_1 ( .OUT(na1884_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3182_1),
                      .CINX(1'b0), .CINY1(na1882_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1884_4 ( .OUT(na1884_2), .IN1(1'b1), .IN2(na3181_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3182_1),
                      .CINX(1'b0), .CINY1(na1882_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x89y71     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1885_2 ( .OUT(na1885_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1885_6 ( .COUTY1(na1885_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1885_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x95y69     80'h00_0078_00_0020_0C66_AAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1886_1 ( .OUT(na1886_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4385_2), .IN6(1'b1), .IN7(na3170_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1888_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1886_4 ( .OUT(na1886_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3172_2), .IN5(na4385_2), .IN6(1'b1), .IN7(na3170_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1888_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x95y68     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1888_2 ( .OUT(na1888_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1888_6 ( .COUTY1(na1888_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1888_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x143y69     80'h00_0078_00_0020_0C66_AC0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1890_1 ( .OUT(na1890_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3213_1), .IN7(na3212_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1899_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1890_4 ( .OUT(na1890_2), .COUTY1(na1890_4), .IN1(na3214_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3213_1),
                      .IN7(na3212_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1899_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y70     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1892_1 ( .OUT(na1892_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3215_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1890_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1892_4 ( .OUT(na1892_2), .COUTY1(na1892_4), .IN1(1'b0), .IN2(1'b0), .IN3(na3216_1), .IN4(1'b1), .IN5(na3215_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1890_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y71     80'h00_0078_00_0020_0C66_0C0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1894_1 ( .OUT(na1894_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3217_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1892_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1894_4 ( .OUT(na1894_2), .COUTY1(na1894_4), .IN1(na3214_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3217_1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1892_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y72     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1896_1 ( .OUT(na1896_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3219_2),
                      .CINX(1'b0), .CINY1(na1894_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1896_4 ( .OUT(na1896_2), .COUTY1(na1896_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3220_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na3219_2), .CINX(1'b0), .CINY1(na1894_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y73     80'h00_0078_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1898_1 ( .OUT(na1898_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3220_2),
                      .CINX(1'b0), .CINY1(na1896_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1898_4 ( .OUT(na1898_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3216_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3220_2),
                      .CINX(1'b0), .CINY1(na1896_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x143y68     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1899_2 ( .OUT(na1899_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1899_6 ( .COUTY1(na1899_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1899_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x144y76     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1900_1 ( .OUT(na1900_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3235_2), .IN6(1'b1), .IN7(1'b1), .IN8(na4393_2),
                      .CINX(1'b0), .CINY1(na3280_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1900_4 ( .OUT(na1900_2), .IN1(na3235_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3235_2), .IN6(1'b1), .IN7(1'b1), .IN8(na4393_2),
                      .CINX(1'b0), .CINY1(na3280_4), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x103y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1903_4 ( .OUT(na1903_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1903_5 ( .OUT(na1903_2), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1903_2_i) );
// C_AND/D///      x126y102     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1904_1 ( .OUT(na1904_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1904_2 ( .OUT(na1904_1), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1904_1_i) );
// C_///AND/D      x108y106     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1905_4 ( .OUT(na1905_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1905_5 ( .OUT(na1905_2), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1905_2_i) );
// C_AND/D///      x101y109     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1906_1 ( .OUT(na1906_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1906_2 ( .OUT(na1906_1), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1906_1_i) );
// C_///AND/D      x98y90     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1907_4 ( .OUT(na1907_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1907_5 ( .OUT(na1907_2), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1907_2_i) );
// C_AND/D///      x97y72     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1908_1 ( .OUT(na1908_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1908_2 ( .OUT(na1908_1), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1908_1_i) );
// C_///AND/D      x101y86     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1909_4 ( .OUT(na1909_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1909_5 ( .OUT(na1909_2), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1909_2_i) );
// C_AND/D///      x91y77     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1910_1 ( .OUT(na1910_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1910_2 ( .OUT(na1910_1), .CLK(1'b0), .EN(na1375_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1910_1_i) );
// C_///AND/D      x149y92     80'h40_F800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1911_4 ( .OUT(na1911_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1134_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1911_5 ( .OUT(na1911_2), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1911_2_i) );
// C_AND/D///      x97y110     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1912_1 ( .OUT(na1912_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1912_2 ( .OUT(na1912_1), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1912_1_i) );
// C_///AND/D      x127y106     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1913_4 ( .OUT(na1913_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1913_5 ( .OUT(na1913_2), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1913_2_i) );
// C_AND/D///      x113y111     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1914_1 ( .OUT(na1914_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1914_2 ( .OUT(na1914_1), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1914_1_i) );
// C_///AND/D      x97y110     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1915_4 ( .OUT(na1915_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1915_5 ( .OUT(na1915_2), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1915_2_i) );
// C_AND/D///      x97y93     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1916_1 ( .OUT(na1916_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1916_2 ( .OUT(na1916_1), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1916_1_i) );
// C_///AND/D      x99y73     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1917_4 ( .OUT(na1917_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1917_5 ( .OUT(na1917_2), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1917_2_i) );
// C_AND/D///      x95y92     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1918_1 ( .OUT(na1918_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1918_2 ( .OUT(na1918_1), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1918_1_i) );
// C_///AND/D      x91y70     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1919_4 ( .OUT(na1919_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1919_5 ( .OUT(na1919_2), .CLK(1'b0), .EN(na1467_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1919_2_i) );
// C_AND/D///      x135y90     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1920_1 ( .OUT(na1920_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1093_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1920_2 ( .OUT(na1920_1), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1920_1_i) );
// C_///AND/D      x141y91     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1921_4 ( .OUT(na1921_2_i), .IN1(1'b1), .IN2(na1094_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1921_5 ( .OUT(na1921_2), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1921_2_i) );
// C_AND/D///      x139y84     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1922_1 ( .OUT(na1922_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1095_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1922_2 ( .OUT(na1922_1), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1922_1_i) );
// C_///AND/D      x136y88     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1923_4 ( .OUT(na1923_2_i), .IN1(1'b1), .IN2(na1096_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1923_5 ( .OUT(na1923_2), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1923_2_i) );
// C_AND/D///      x139y76     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1924_1 ( .OUT(na1924_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1097_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1924_2 ( .OUT(na1924_1), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1924_1_i) );
// C_///AND/D      x138y70     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1925_4 ( .OUT(na1925_2_i), .IN1(na1098_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1925_5 ( .OUT(na1925_2), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1925_2_i) );
// C_AND/D///      x137y83     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1926_1 ( .OUT(na1926_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1099_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1926_2 ( .OUT(na1926_1), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1926_1_i) );
// C_///AND/D      x136y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1927_4 ( .OUT(na1927_2_i), .IN1(1'b1), .IN2(na1100_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1927_5 ( .OUT(na1927_2), .CLK(1'b0), .EN(na1456_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1927_2_i) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0000_0010)) 
           _a1928 ( .GLB0(na1928_1), .GLB1(_d3), .GLB2(_d4), .GLB3(_d5), .CLK_FB0(_d6), .CLK_FB1(_d7), .CLK_FB2(_d8), .CLK_FB3(_d9),
                    .CLK0_0(1'b0), .CLK0_90(1'b0), .CLK0_180(1'b0), .CLK0_270(1'b0), .CLK0_BYP(na14_1), .CLK1_0(1'b0), .CLK1_90(1'b0),
                    .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                    .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(1'b0),
                    .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_AND/D///      x149y82     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1929_1 ( .OUT(na1929_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1929_2 ( .OUT(na1929_1), .CLK(1'b0), .EN(na1455_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1929_1_i) );
// C_AND/D//AND/D      x148y81     80'h40_E800_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1930_1 ( .OUT(na1930_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1930_2 ( .OUT(na1930_1), .CLK(1'b0), .EN(na1455_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1930_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1930_4 ( .OUT(na1930_2_i), .IN1(1'b1), .IN2(na8_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1930_5 ( .OUT(na1930_2), .CLK(1'b0), .EN(na1455_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1930_2_i) );
// C_AND/D//AND/D      x148y84     80'h40_E800_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1932_1 ( .OUT(na1932_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na12_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1932_2 ( .OUT(na1932_1), .CLK(1'b0), .EN(na1455_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1932_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1932_4 ( .OUT(na1932_2_i), .IN1(na11_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1932_5 ( .OUT(na1932_2), .CLK(1'b0), .EN(na1455_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1932_2_i) );
// C_///AND/D      x92y98     80'h40_E400_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1934_4 ( .OUT(na1934_2_i), .IN1(1'b1), .IN2(na2_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1934_5 ( .OUT(na1934_2), .CLK(1'b0), .EN(~na1454_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1934_2_i) );
// C_AND/D//AND/D      x89y103     80'h40_E400_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1935_1 ( .OUT(na1935_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1935_2 ( .OUT(na1935_1), .CLK(1'b0), .EN(~na1454_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1935_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1935_4 ( .OUT(na1935_2_i), .IN1(1'b1), .IN2(na1_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1935_5 ( .OUT(na1935_2), .CLK(1'b0), .EN(~na1454_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1935_2_i) );
// C_AND/D//AND/D      x91y106     80'h40_E400_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1937_1 ( .OUT(na1937_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1937_2 ( .OUT(na1937_1), .CLK(1'b0), .EN(~na1454_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1937_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1937_4 ( .OUT(na1937_2_i), .IN1(1'b1), .IN2(na4_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1937_5 ( .OUT(na1937_2), .CLK(1'b0), .EN(~na1454_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1937_2_i) );
// C_AND/D///      x92y110     80'h40_E400_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1938_1 ( .OUT(na1938_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1938_2 ( .OUT(na1938_1), .CLK(1'b0), .EN(~na1454_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1938_1_i) );
// C_AND/D//AND/D      x149y96     80'h40_E800_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1941_1 ( .OUT(na1941_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1248_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1941_2 ( .OUT(na1941_1), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1941_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1941_4 ( .OUT(na1941_2_i), .IN1(1'b1), .IN2(na1203_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1941_5 ( .OUT(na1941_2), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1941_2_i) );
// C_AND/D//AND/D      x146y95     80'h40_E800_80_0000_0C88_F3FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1943_1 ( .OUT(na1943_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1271_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1943_2 ( .OUT(na1943_1), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1943_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1943_4 ( .OUT(na1943_2_i), .IN1(1'b1), .IN2(na1260_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1943_5 ( .OUT(na1943_2), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1943_2_i) );
// C_AND/D//AND/D      x145y95     80'h40_E800_80_0000_0C88_FA3F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1945_1 ( .OUT(na1945_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1293_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1945_2 ( .OUT(na1945_1), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1945_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1945_4 ( .OUT(na1945_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1282_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1945_5 ( .OUT(na1945_2), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1945_2_i) );
// C_AND/D//AND/D      x144y96     80'h40_E800_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1946_1 ( .OUT(na1946_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1304_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1946_2 ( .OUT(na1946_1), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1946_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1946_4 ( .OUT(na1946_2_i), .IN1(na1237_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1946_5 ( .OUT(na1946_2), .CLK(1'b0), .EN(na7_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1946_2_i) );
// C_///AND/D      x148y69     80'h40_E800_80_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1947_4 ( .OUT(na1947_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1374_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1947_5 ( .OUT(na1947_2), .CLK(1'b0), .EN(na1958_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1947_2_i) );
// C_AND/D///      x120y76     80'h40_E400_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1948_1 ( .OUT(na1948_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1373_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1948_2 ( .OUT(na1948_1), .CLK(1'b0), .EN(~na1457_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1948_1_i) );
// C_///AND/D      x112y101     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1949_4 ( .OUT(na1949_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1949_5 ( .OUT(na1949_2), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1949_2_i) );
// C_AND/D///      x122y99     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1950_1 ( .OUT(na1950_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1950_2 ( .OUT(na1950_1), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1950_1_i) );
// C_///AND/D      x91y103     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1951_4 ( .OUT(na1951_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1951_5 ( .OUT(na1951_2), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1951_2_i) );
// C_AND/D///      x102y106     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1952_1 ( .OUT(na1952_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1952_2 ( .OUT(na1952_1), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1952_1_i) );
// C_///AND/D      x105y99     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1953_4 ( .OUT(na1953_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1953_5 ( .OUT(na1953_2), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1953_2_i) );
// C_AND/D///      x100y72     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1954_1 ( .OUT(na1954_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1954_2 ( .OUT(na1954_1), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1954_1_i) );
// C_///AND/D      x105y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1955_4 ( .OUT(na1955_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1955_5 ( .OUT(na1955_2), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1955_2_i) );
// C_AND/D///      x94y80     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1956_1 ( .OUT(na1956_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1956_2 ( .OUT(na1956_1), .CLK(1'b0), .EN(na1409_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1956_1_i) );
// C_///AND/D      x139y66     80'h40_EC00_80_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1957_4 ( .OUT(na1957_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na531_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1957_5 ( .OUT(na1957_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1957_2_i) );
// C_AND/D///      x142y67     80'h40_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1958_1 ( .OUT(na1958_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na540_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1958_2 ( .OUT(na1958_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1958_1_i) );
// C_///AND/D      x100y102     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1959_4 ( .OUT(na1959_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1959_5 ( .OUT(na1959_2), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1959_2_i) );
// C_AND/D///      x122y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1960_1 ( .OUT(na1960_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1960_2 ( .OUT(na1960_1), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1960_1_i) );
// C_///AND/D      x106y102     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1961_4 ( .OUT(na1961_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1961_5 ( .OUT(na1961_2), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1961_2_i) );
// C_AND/D///      x100y102     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1962_1 ( .OUT(na1962_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1962_2 ( .OUT(na1962_1), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1962_1_i) );
// C_///AND/D      x100y82     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1963_4 ( .OUT(na1963_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1963_5 ( .OUT(na1963_2), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1963_2_i) );
// C_AND/D///      x100y74     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1964_1 ( .OUT(na1964_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1964_2 ( .OUT(na1964_1), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1964_1_i) );
// C_///AND/D      x100y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1965_4 ( .OUT(na1965_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1965_5 ( .OUT(na1965_2), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1965_2_i) );
// C_AND/D///      x96y72     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1966_1 ( .OUT(na1966_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1966_2 ( .OUT(na1966_1), .CLK(1'b0), .EN(na1390_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1966_1_i) );
// C_///AND/D      x96y104     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1967_4 ( .OUT(na1967_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1967_5 ( .OUT(na1967_2), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1967_2_i) );
// C_AND/D///      x118y102     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1968_1 ( .OUT(na1968_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1968_2 ( .OUT(na1968_1), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1968_1_i) );
// C_///AND/D      x108y98     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1969_4 ( .OUT(na1969_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1969_5 ( .OUT(na1969_2), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1969_2_i) );
// C_AND/D///      x97y102     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1970_1 ( .OUT(na1970_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1970_2 ( .OUT(na1970_1), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1970_1_i) );
// C_///AND/D      x98y80     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1971_4 ( .OUT(na1971_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1971_5 ( .OUT(na1971_2), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1971_2_i) );
// C_AND/D///      x98y76     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1972_1 ( .OUT(na1972_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1972_2 ( .OUT(na1972_1), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1972_1_i) );
// C_///AND/D      x104y80     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1973_4 ( .OUT(na1973_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1973_5 ( .OUT(na1973_2), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1973_2_i) );
// C_AND/D///      x96y78     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1974_1 ( .OUT(na1974_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1974_2 ( .OUT(na1974_1), .CLK(1'b0), .EN(na1391_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1974_1_i) );
// C_///AND/D      x93y101     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1975_4 ( .OUT(na1975_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1975_5 ( .OUT(na1975_2), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1975_2_i) );
// C_AND/D///      x113y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1976_1 ( .OUT(na1976_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1976_2 ( .OUT(na1976_1), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1976_1_i) );
// C_///AND/D      x103y101     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1977_4 ( .OUT(na1977_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1977_5 ( .OUT(na1977_2), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1977_2_i) );
// C_AND/D///      x102y100     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1978_1 ( .OUT(na1978_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1978_2 ( .OUT(na1978_1), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1978_1_i) );
// C_///AND/D      x87y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1979_4 ( .OUT(na1979_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1979_5 ( .OUT(na1979_2), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1979_2_i) );
// C_AND/D///      x102y72     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1980_1 ( .OUT(na1980_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1980_2 ( .OUT(na1980_1), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1980_1_i) );
// C_///AND/D      x93y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1981_4 ( .OUT(na1981_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1981_5 ( .OUT(na1981_2), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1981_2_i) );
// C_AND/D///      x87y72     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1982_1 ( .OUT(na1982_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1982_2 ( .OUT(na1982_1), .CLK(1'b0), .EN(na1393_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1982_1_i) );
// C_///AND/D      x102y103     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1983_4 ( .OUT(na1983_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1983_5 ( .OUT(na1983_2), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1983_2_i) );
// C_AND/D///      x120y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1984_1 ( .OUT(na1984_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1984_2 ( .OUT(na1984_1), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1984_1_i) );
// C_///AND/D      x108y99     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1985_4 ( .OUT(na1985_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1985_5 ( .OUT(na1985_2), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1985_2_i) );
// C_AND/D///      x102y103     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1986_1 ( .OUT(na1986_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1986_2 ( .OUT(na1986_1), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1986_1_i) );
// C_///AND/D      x96y87     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1987_4 ( .OUT(na1987_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1987_5 ( .OUT(na1987_2), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1987_2_i) );
// C_AND/D///      x100y77     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1988_1 ( .OUT(na1988_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1988_2 ( .OUT(na1988_1), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1988_1_i) );
// C_///AND/D      x98y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1989_4 ( .OUT(na1989_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1989_5 ( .OUT(na1989_2), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1989_2_i) );
// C_AND/D///      x96y77     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1990_1 ( .OUT(na1990_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1990_2 ( .OUT(na1990_1), .CLK(1'b0), .EN(na1394_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1990_1_i) );
// C_AND/D///      x100y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1991_1 ( .OUT(na1991_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1991_2 ( .OUT(na1991_1), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1991_1_i) );
// C_AND/D///      x118y103     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1992_1 ( .OUT(na1992_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1992_2 ( .OUT(na1992_1), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1992_1_i) );
// C_///AND/D      x104y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1993_4 ( .OUT(na1993_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1993_5 ( .OUT(na1993_2), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1993_2_i) );
// C_AND/D///      x98y101     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1994_1 ( .OUT(na1994_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1994_2 ( .OUT(na1994_1), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1994_1_i) );
// C_///AND/D      x98y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1995_4 ( .OUT(na1995_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1995_5 ( .OUT(na1995_2), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1995_2_i) );
// C_AND/D///      x100y73     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1996_1 ( .OUT(na1996_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1996_2 ( .OUT(na1996_1), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1996_1_i) );
// C_///AND/D      x100y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1997_4 ( .OUT(na1997_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1997_5 ( .OUT(na1997_2), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1997_2_i) );
// C_AND/D///      x94y73     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1998_1 ( .OUT(na1998_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1998_2 ( .OUT(na1998_1), .CLK(1'b0), .EN(na1396_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1998_1_i) );
// C_///AND/D      x102y101     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1999_4 ( .OUT(na1999_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1999_5 ( .OUT(na1999_2), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1999_2_i) );
// C_AND/D///      x122y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2000_1 ( .OUT(na2000_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2000_2 ( .OUT(na2000_1), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2000_1_i) );
// C_///AND/D      x106y99     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2001_4 ( .OUT(na2001_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2001_5 ( .OUT(na2001_2), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2001_2_i) );
// C_AND/D///      x98y103     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2002_1 ( .OUT(na2002_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2002_2 ( .OUT(na2002_1), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2002_1_i) );
// C_///AND/D      x96y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2003_4 ( .OUT(na2003_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2003_5 ( .OUT(na2003_2), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2003_2_i) );
// C_AND/D///      x98y75     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2004_1 ( .OUT(na2004_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2004_2 ( .OUT(na2004_1), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2004_1_i) );
// C_///AND/D      x102y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2005_4 ( .OUT(na2005_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2005_5 ( .OUT(na2005_2), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2005_2_i) );
// C_AND/D///      x92y73     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2006_1 ( .OUT(na2006_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2006_2 ( .OUT(na2006_1), .CLK(1'b0), .EN(na1397_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2006_1_i) );
// C_///AND/D      x94y101     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2007_4 ( .OUT(na2007_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2007_5 ( .OUT(na2007_2), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2007_2_i) );
// C_AND/D///      x114y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2008_1 ( .OUT(na2008_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2008_2 ( .OUT(na2008_1), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2008_1_i) );
// C_///AND/D      x104y95     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2009_4 ( .OUT(na2009_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2009_5 ( .OUT(na2009_2), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2009_2_i) );
// C_AND/D///      x94y103     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2010_1 ( .OUT(na2010_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2010_2 ( .OUT(na2010_1), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2010_1_i) );
// C_///AND/D      x94y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2011_4 ( .OUT(na2011_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2011_5 ( .OUT(na2011_2), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2011_2_i) );
// C_AND/D///      x102y81     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2012_1 ( .OUT(na2012_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2012_2 ( .OUT(na2012_1), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2012_1_i) );
// C_///AND/D      x96y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2013_4 ( .OUT(na2013_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2013_5 ( .OUT(na2013_2), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2013_2_i) );
// C_AND/D///      x100y81     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2014_1 ( .OUT(na2014_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2014_2 ( .OUT(na2014_1), .CLK(1'b0), .EN(na1398_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2014_1_i) );
// C_///AND/D      x97y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2015_4 ( .OUT(na2015_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2015_5 ( .OUT(na2015_2), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2015_2_i) );
// C_AND/D///      x117y99     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2016_1 ( .OUT(na2016_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2016_2 ( .OUT(na2016_1), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2016_1_i) );
// C_///AND/D      x111y99     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2017_4 ( .OUT(na2017_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2017_5 ( .OUT(na2017_2), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2017_2_i) );
// C_AND/D///      x100y104     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2018_1 ( .OUT(na2018_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2018_2 ( .OUT(na2018_1), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2018_1_i) );
// C_///AND/D      x99y89     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2019_4 ( .OUT(na2019_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2019_5 ( .OUT(na2019_2), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2019_2_i) );
// C_AND/D///      x97y77     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2020_1 ( .OUT(na2020_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2020_2 ( .OUT(na2020_1), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2020_1_i) );
// C_///AND/D      x99y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2021_4 ( .OUT(na2021_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2021_5 ( .OUT(na2021_2), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2021_2_i) );
// C_AND/D///      x95y77     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2022_1 ( .OUT(na2022_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2022_2 ( .OUT(na2022_1), .CLK(1'b0), .EN(na1399_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2022_1_i) );
// C_///AND/D      x103y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2023_4 ( .OUT(na2023_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2023_5 ( .OUT(na2023_2), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2023_2_i) );
// C_AND/D///      x119y103     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2024_1 ( .OUT(na2024_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2024_2 ( .OUT(na2024_1), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2024_1_i) );
// C_///AND/D      x105y101     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2025_4 ( .OUT(na2025_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2025_5 ( .OUT(na2025_2), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2025_2_i) );
// C_AND/D///      x99y103     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2026_1 ( .OUT(na2026_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2026_2 ( .OUT(na2026_1), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2026_1_i) );
// C_///AND/D      x97y83     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2027_4 ( .OUT(na2027_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2027_5 ( .OUT(na2027_2), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2027_2_i) );
// C_AND/D///      x101y73     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2028_1 ( .OUT(na2028_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2028_2 ( .OUT(na2028_1), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2028_1_i) );
// C_///AND/D      x101y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2029_4 ( .OUT(na2029_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2029_5 ( .OUT(na2029_2), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2029_2_i) );
// C_AND/D///      x95y73     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2030_1 ( .OUT(na2030_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2030_2 ( .OUT(na2030_1), .CLK(1'b0), .EN(na1401_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2030_1_i) );
// C_///AND/D      x99y105     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2031_4 ( .OUT(na2031_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2031_5 ( .OUT(na2031_2), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2031_2_i) );
// C_AND/D///      x121y103     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2032_1 ( .OUT(na2032_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2032_2 ( .OUT(na2032_1), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2032_1_i) );
// C_///AND/D      x107y105     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2033_4 ( .OUT(na2033_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2033_5 ( .OUT(na2033_2), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2033_2_i) );
// C_AND/D///      x98y104     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2034_1 ( .OUT(na2034_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2034_2 ( .OUT(na2034_1), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2034_1_i) );
// C_///AND/D      x95y81     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2035_4 ( .OUT(na2035_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2035_5 ( .OUT(na2035_2), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2035_2_i) );
// C_AND/D///      x101y75     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2036_1 ( .OUT(na2036_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2036_2 ( .OUT(na2036_1), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2036_1_i) );
// C_///AND/D      x103y77     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2037_4 ( .OUT(na2037_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2037_5 ( .OUT(na2037_2), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2037_2_i) );
// C_AND/D///      x93y75     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2038_1 ( .OUT(na2038_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2038_2 ( .OUT(na2038_1), .CLK(1'b0), .EN(na1402_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2038_1_i) );
// C_///AND/D      x97y103     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2039_4 ( .OUT(na2039_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2039_5 ( .OUT(na2039_2), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2039_2_i) );
// C_AND/D///      x119y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2040_1 ( .OUT(na2040_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2040_2 ( .OUT(na2040_1), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2040_1_i) );
// C_///AND/D      x101y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2041_4 ( .OUT(na2041_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2041_5 ( .OUT(na2041_2), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2041_2_i) );
// C_AND/D///      x95y105     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2042_1 ( .OUT(na2042_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2042_2 ( .OUT(na2042_1), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2042_1_i) );
// C_///AND/D      x89y81     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2043_4 ( .OUT(na2043_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2043_5 ( .OUT(na2043_2), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2043_2_i) );
// C_AND/D///      x99y77     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2044_1 ( .OUT(na2044_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2044_2 ( .OUT(na2044_1), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2044_1_i) );
// C_///AND/D      x95y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2045_4 ( .OUT(na2045_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2045_5 ( .OUT(na2045_2), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2045_2_i) );
// C_AND/D///      x97y79     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2046_1 ( .OUT(na2046_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2046_2 ( .OUT(na2046_1), .CLK(1'b0), .EN(na1403_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2046_1_i) );
// C_///AND/D      x99y100     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2047_4 ( .OUT(na2047_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2047_5 ( .OUT(na2047_2), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2047_2_i) );
// C_AND/D///      x117y100     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2048_1 ( .OUT(na2048_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2048_2 ( .OUT(na2048_1), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2048_1_i) );
// C_///AND/D      x107y96     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2049_4 ( .OUT(na2049_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2049_5 ( .OUT(na2049_2), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2049_2_i) );
// C_AND/D///      x99y104     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2050_1 ( .OUT(na2050_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2050_2 ( .OUT(na2050_1), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2050_1_i) );
// C_///AND/D      x99y86     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2051_4 ( .OUT(na2051_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2051_5 ( .OUT(na2051_2), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2051_2_i) );
// C_AND/D///      x99y76     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2052_1 ( .OUT(na2052_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2052_2 ( .OUT(na2052_1), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2052_1_i) );
// C_///AND/D      x101y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2053_4 ( .OUT(na2053_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2053_5 ( .OUT(na2053_2), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2053_2_i) );
// C_AND/D///      x93y78     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2054_1 ( .OUT(na2054_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2054_2 ( .OUT(na2054_1), .CLK(1'b0), .EN(na1404_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2054_1_i) );
// C_///AND/D      x99y102     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2055_4 ( .OUT(na2055_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2055_5 ( .OUT(na2055_2), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2055_2_i) );
// C_AND/D///      x117y102     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2056_1 ( .OUT(na2056_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2056_2 ( .OUT(na2056_1), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2056_1_i) );
// C_///AND/D      x105y102     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2057_4 ( .OUT(na2057_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2057_5 ( .OUT(na2057_2), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2057_2_i) );
// C_AND/D///      x97y104     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2058_1 ( .OUT(na2058_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2058_2 ( .OUT(na2058_1), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2058_1_i) );
// C_///AND/D      x101y84     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2059_4 ( .OUT(na2059_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2059_5 ( .OUT(na2059_2), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2059_2_i) );
// C_AND/D///      x99y74     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2060_1 ( .OUT(na2060_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2060_2 ( .OUT(na2060_1), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2060_1_i) );
// C_///AND/D      x95y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2061_4 ( .OUT(na2061_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2061_5 ( .OUT(na2061_2), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2061_2_i) );
// C_AND/D///      x95y74     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2062_1 ( .OUT(na2062_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2062_2 ( .OUT(na2062_1), .CLK(1'b0), .EN(na1412_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2062_1_i) );
// C_///AND/D      x85y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2063_4 ( .OUT(na2063_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2063_5 ( .OUT(na2063_2), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2063_2_i) );
// C_AND/D///      x122y112     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2064_1 ( .OUT(na2064_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2064_2 ( .OUT(na2064_1), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2064_1_i) );
// C_///AND/D      x104y109     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2065_4 ( .OUT(na2065_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2065_5 ( .OUT(na2065_2), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2065_2_i) );
// C_AND/D///      x97y113     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2066_1 ( .OUT(na2066_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2066_2 ( .OUT(na2066_1), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2066_1_i) );
// C_///AND/D      x92y102     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2067_4 ( .OUT(na2067_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2067_5 ( .OUT(na2067_2), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2067_2_i) );
// C_AND/D///      x89y84     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2068_1 ( .OUT(na2068_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2068_2 ( .OUT(na2068_1), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2068_1_i) );
// C_///AND/D      x90y90     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2069_4 ( .OUT(na2069_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2069_5 ( .OUT(na2069_2), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2069_2_i) );
// C_AND/D///      x87y83     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2070_1 ( .OUT(na2070_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2070_2 ( .OUT(na2070_1), .CLK(1'b0), .EN(na1405_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2070_1_i) );
// C_///AND/D      x90y102     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2071_4 ( .OUT(na2071_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2071_5 ( .OUT(na2071_2), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2071_2_i) );
// C_AND/D///      x107y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2072_1 ( .OUT(na2072_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2072_2 ( .OUT(na2072_1), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2072_1_i) );
// C_///AND/D      x98y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2073_4 ( .OUT(na2073_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2073_5 ( .OUT(na2073_2), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2073_2_i) );
// C_AND/D///      x93y105     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2074_1 ( .OUT(na2074_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2074_2 ( .OUT(na2074_1), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2074_1_i) );
// C_///AND/D      x88y82     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2075_4 ( .OUT(na2075_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2075_5 ( .OUT(na2075_2), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2075_2_i) );
// C_AND/D///      x97y78     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2076_1 ( .OUT(na2076_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2076_2 ( .OUT(na2076_1), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2076_1_i) );
// C_///AND/D      x90y83     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2077_4 ( .OUT(na2077_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2077_5 ( .OUT(na2077_2), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2077_2_i) );
// C_AND/D///      x97y69     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2078_1 ( .OUT(na2078_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2078_2 ( .OUT(na2078_1), .CLK(1'b0), .EN(na1407_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2078_1_i) );
// C_///AND/D      x100y106     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2079_4 ( .OUT(na2079_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2079_5 ( .OUT(na2079_2), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2079_2_i) );
// C_AND/D///      x120y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2080_1 ( .OUT(na2080_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2080_2 ( .OUT(na2080_1), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2080_1_i) );
// C_///AND/D      x114y109     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2081_4 ( .OUT(na2081_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2081_5 ( .OUT(na2081_2), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2081_2_i) );
// C_AND/D///      x99y106     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2082_1 ( .OUT(na2082_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2082_2 ( .OUT(na2082_1), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2082_1_i) );
// C_///AND/D      x106y91     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2083_4 ( .OUT(na2083_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2083_5 ( .OUT(na2083_2), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2083_2_i) );
// C_AND/D///      x100y80     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2084_1 ( .OUT(na2084_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2084_2 ( .OUT(na2084_1), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2084_1_i) );
// C_///AND/D      x104y91     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2085_4 ( .OUT(na2085_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2085_5 ( .OUT(na2085_2), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2085_2_i) );
// C_AND/D///      x92y76     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2086_1 ( .OUT(na2086_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2086_2 ( .OUT(na2086_1), .CLK(1'b0), .EN(na1408_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2086_1_i) );
// C_///AND/D      x98y95     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2087_4 ( .OUT(na2087_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2087_5 ( .OUT(na2087_2), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2087_2_i) );
// C_AND/D///      x119y94     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2088_1 ( .OUT(na2088_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2088_2 ( .OUT(na2088_1), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2088_1_i) );
// C_///AND/D      x102y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2089_4 ( .OUT(na2089_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2089_5 ( .OUT(na2089_2), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2089_2_i) );
// C_AND/D///      x94y102     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2090_1 ( .OUT(na2090_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2090_2 ( .OUT(na2090_1), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2090_1_i) );
// C_///AND/D      x102y78     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2091_4 ( .OUT(na2091_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2091_5 ( .OUT(na2091_2), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2091_2_i) );
// C_AND/D///      x97y67     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2092_1 ( .OUT(na2092_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2092_2 ( .OUT(na2092_1), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2092_1_i) );
// C_///AND/D      x96y83     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2093_4 ( .OUT(na2093_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2093_5 ( .OUT(na2093_2), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2093_2_i) );
// C_AND/D///      x92y69     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2094_1 ( .OUT(na2094_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2094_2 ( .OUT(na2094_1), .CLK(1'b0), .EN(na1410_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2094_1_i) );
// C_///AND/D      x101y106     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2095_4 ( .OUT(na2095_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2095_5 ( .OUT(na2095_2), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2095_2_i) );
// C_AND/D///      x119y102     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2096_1 ( .OUT(na2096_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2096_2 ( .OUT(na2096_1), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2096_1_i) );
// C_///AND/D      x107y104     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2097_4 ( .OUT(na2097_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2097_5 ( .OUT(na2097_2), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2097_2_i) );
// C_AND/D///      x95y102     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2098_1 ( .OUT(na2098_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2098_2 ( .OUT(na2098_1), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2098_1_i) );
// C_///AND/D      x97y82     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2099_4 ( .OUT(na2099_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2099_5 ( .OUT(na2099_2), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2099_2_i) );
// C_AND/D///      x103y78     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2100_1 ( .OUT(na2100_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2100_2 ( .OUT(na2100_1), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2100_1_i) );
// C_///AND/D      x103y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2101_4 ( .OUT(na2101_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2101_5 ( .OUT(na2101_2), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2101_2_i) );
// C_AND/D///      x97y74     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2102_1 ( .OUT(na2102_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2102_2 ( .OUT(na2102_1), .CLK(1'b0), .EN(na1411_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2102_1_i) );
// C_///AND/D      x111y108     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2103_4 ( .OUT(na2103_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2103_5 ( .OUT(na2103_2), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2103_2_i) );
// C_AND/D///      x123y103     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2104_1 ( .OUT(na2104_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2104_2 ( .OUT(na2104_1), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2104_1_i) );
// C_///AND/D      x109y109     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2105_4 ( .OUT(na2105_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2105_5 ( .OUT(na2105_2), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2105_2_i) );
// C_AND/D///      x97y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2106_1 ( .OUT(na2106_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2106_2 ( .OUT(na2106_1), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2106_1_i) );
// C_///AND/D      x103y91     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2107_4 ( .OUT(na2107_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2107_5 ( .OUT(na2107_2), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2107_2_i) );
// C_AND/D///      x99y70     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2108_1 ( .OUT(na2108_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2108_2 ( .OUT(na2108_1), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2108_1_i) );
// C_///AND/D      x103y80     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2109_4 ( .OUT(na2109_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2109_5 ( .OUT(na2109_2), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2109_2_i) );
// C_AND/D///      x87y77     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2110_1 ( .OUT(na2110_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2110_2 ( .OUT(na2110_1), .CLK(1'b0), .EN(na1413_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2110_1_i) );
// C_///AND/D      x89y106     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2111_4 ( .OUT(na2111_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2111_5 ( .OUT(na2111_2), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2111_2_i) );
// C_AND/D///      x107y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2112_1 ( .OUT(na2112_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2112_2 ( .OUT(na2112_1), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2112_1_i) );
// C_///AND/D      x100y93     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2113_4 ( .OUT(na2113_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2113_5 ( .OUT(na2113_2), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2113_2_i) );
// C_AND/D///      x91y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2114_1 ( .OUT(na2114_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2114_2 ( .OUT(na2114_1), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2114_1_i) );
// C_///AND/D      x93y83     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2115_4 ( .OUT(na2115_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2115_5 ( .OUT(na2115_2), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2115_2_i) );
// C_AND/D///      x90y80     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2116_1 ( .OUT(na2116_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2116_2 ( .OUT(na2116_1), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2116_1_i) );
// C_///AND/D      x87y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2117_4 ( .OUT(na2117_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2117_5 ( .OUT(na2117_2), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2117_2_i) );
// C_AND/D///      x87y78     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2118_1 ( .OUT(na2118_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2118_2 ( .OUT(na2118_1), .CLK(1'b0), .EN(na1414_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2118_1_i) );
// C_///AND/D      x101y115     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2119_4 ( .OUT(na2119_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2119_5 ( .OUT(na2119_2), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2119_2_i) );
// C_AND/D///      x125y105     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2120_1 ( .OUT(na2120_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2120_2 ( .OUT(na2120_1), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2120_1_i) );
// C_///AND/D      x113y103     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2121_4 ( .OUT(na2121_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2121_5 ( .OUT(na2121_2), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2121_2_i) );
// C_AND/D///      x95y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2122_1 ( .OUT(na2122_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2122_2 ( .OUT(na2122_1), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2122_1_i) );
// C_///AND/D      x102y94     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2123_4 ( .OUT(na2123_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2123_5 ( .OUT(na2123_2), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2123_2_i) );
// C_AND/D///      x97y76     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2124_1 ( .OUT(na2124_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2124_2 ( .OUT(na2124_1), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2124_1_i) );
// C_///AND/D      x105y94     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2125_4 ( .OUT(na2125_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2125_5 ( .OUT(na2125_2), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2125_2_i) );
// C_AND/D///      x90y78     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2126_1 ( .OUT(na2126_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2126_2 ( .OUT(na2126_1), .CLK(1'b0), .EN(na1415_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2126_1_i) );
// C_///AND/D      x108y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2127_4 ( .OUT(na2127_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2127_5 ( .OUT(na2127_2), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2127_2_i) );
// C_AND/D///      x125y102     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2128_1 ( .OUT(na2128_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2128_2 ( .OUT(na2128_1), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2128_1_i) );
// C_///AND/D      x113y106     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2129_4 ( .OUT(na2129_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2129_5 ( .OUT(na2129_2), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2129_2_i) );
// C_AND/D///      x100y111     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2130_1 ( .OUT(na2130_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2130_2 ( .OUT(na2130_1), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2130_1_i) );
// C_///AND/D      x91y88     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2131_4 ( .OUT(na2131_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2131_5 ( .OUT(na2131_2), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2131_2_i) );
// C_AND/D///      x97y68     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2132_1 ( .OUT(na2132_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2132_2 ( .OUT(na2132_1), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2132_1_i) );
// C_///AND/D      x103y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2133_4 ( .OUT(na2133_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2133_5 ( .OUT(na2133_2), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2133_2_i) );
// C_AND/D///      x87y80     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2134_1 ( .OUT(na2134_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2134_2 ( .OUT(na2134_1), .CLK(1'b0), .EN(na1416_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2134_1_i) );
// C_///AND/D      x93y112     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2135_4 ( .OUT(na2135_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2135_5 ( .OUT(na2135_2), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2135_2_i) );
// C_///AND/D      x127y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2136_4 ( .OUT(na2136_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2136_5 ( .OUT(na2136_2), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2136_2_i) );
// C_///AND/D      x101y108     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2137_4 ( .OUT(na2137_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2137_5 ( .OUT(na2137_2), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2137_2_i) );
// C_AND/D///      x93y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2138_1 ( .OUT(na2138_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2138_2 ( .OUT(na2138_1), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2138_1_i) );
// C_///AND/D      x95y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2139_4 ( .OUT(na2139_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2139_5 ( .OUT(na2139_2), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2139_2_i) );
// C_AND/D///      x91y82     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2140_1 ( .OUT(na2140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2140_2 ( .OUT(na2140_1), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2140_1_i) );
// C_///AND/D      x88y89     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2141_4 ( .OUT(na2141_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2141_5 ( .OUT(na2141_2), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2141_2_i) );
// C_AND/D///      x85y81     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2142_1 ( .OUT(na2142_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2142_2 ( .OUT(na2142_1), .CLK(1'b0), .EN(na1417_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2142_1_i) );
// C_///AND/D      x89y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2143_4 ( .OUT(na2143_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2143_5 ( .OUT(na2143_2), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2143_2_i) );
// C_AND/D///      x108y108     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2144_1 ( .OUT(na2144_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2144_2 ( .OUT(na2144_1), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2144_1_i) );
// C_///AND/D      x99y94     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2145_4 ( .OUT(na2145_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2145_5 ( .OUT(na2145_2), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2145_2_i) );
// C_AND/D///      x89y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2146_1 ( .OUT(na2146_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2146_2 ( .OUT(na2146_1), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2146_1_i) );
// C_///AND/D      x88y83     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2147_4 ( .OUT(na2147_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2147_5 ( .OUT(na2147_2), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2147_2_i) );
// C_AND/D///      x93y82     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2148_1 ( .OUT(na2148_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2148_2 ( .OUT(na2148_1), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2148_1_i) );
// C_///AND/D      x85y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2149_4 ( .OUT(na2149_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2149_5 ( .OUT(na2149_2), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2149_2_i) );
// C_AND/D///      x91y69     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2150_1 ( .OUT(na2150_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2150_2 ( .OUT(na2150_1), .CLK(1'b0), .EN(na1418_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2150_1_i) );
// C_///AND/D      x101y112     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2151_4 ( .OUT(na2151_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2151_5 ( .OUT(na2151_2), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2151_2_i) );
// C_AND/D///      x123y106     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2152_1 ( .OUT(na2152_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2152_2 ( .OUT(na2152_1), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2152_1_i) );
// C_///AND/D      x114y106     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2153_4 ( .OUT(na2153_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2153_5 ( .OUT(na2153_2), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2153_2_i) );
// C_AND/D///      x101y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2154_1 ( .OUT(na2154_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2154_2 ( .OUT(na2154_1), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2154_1_i) );
// C_///AND/D      x104y94     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2155_4 ( .OUT(na2155_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2155_5 ( .OUT(na2155_2), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2155_2_i) );
// C_AND/D///      x102y77     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2156_1 ( .OUT(na2156_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2156_2 ( .OUT(na2156_1), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2156_1_i) );
// C_///AND/D      x103y89     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2157_4 ( .OUT(na2157_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2157_5 ( .OUT(na2157_2), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2157_2_i) );
// C_AND/D///      x89y80     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2158_1 ( .OUT(na2158_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2158_2 ( .OUT(na2158_1), .CLK(1'b0), .EN(na1419_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2158_1_i) );
// C_///AND/D      x96y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2159_4 ( .OUT(na2159_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2159_5 ( .OUT(na2159_2), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2159_2_i) );
// C_AND/D///      x125y106     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2160_1 ( .OUT(na2160_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2160_2 ( .OUT(na2160_1), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2160_1_i) );
// C_///AND/D      x107y102     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2161_4 ( .OUT(na2161_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2161_5 ( .OUT(na2161_2), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2161_2_i) );
// C_AND/D///      x96y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2162_1 ( .OUT(na2162_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2162_2 ( .OUT(na2162_1), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2162_1_i) );
// C_///AND/D      x96y98     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2163_4 ( .OUT(na2163_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2163_5 ( .OUT(na2163_2), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2163_2_i) );
// C_AND/D///      x94y82     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2164_1 ( .OUT(na2164_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2164_2 ( .OUT(na2164_1), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2164_1_i) );
// C_///AND/D      x91y96     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2165_4 ( .OUT(na2165_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2165_5 ( .OUT(na2165_2), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2165_2_i) );
// C_AND/D///      x90y82     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2166_1 ( .OUT(na2166_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2166_2 ( .OUT(na2166_1), .CLK(1'b0), .EN(na1420_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2166_1_i) );
// C_///AND/D      x100y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2167_4 ( .OUT(na2167_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2167_5 ( .OUT(na2167_2), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2167_2_i) );
// C_AND/D///      x121y106     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2168_1 ( .OUT(na2168_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2168_2 ( .OUT(na2168_1), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2168_1_i) );
// C_///AND/D      x116y106     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2169_4 ( .OUT(na2169_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2169_5 ( .OUT(na2169_2), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2169_2_i) );
// C_AND/D///      x100y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2170_1 ( .OUT(na2170_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2170_2 ( .OUT(na2170_1), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2170_1_i) );
// C_///AND/D      x105y89     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2171_4 ( .OUT(na2171_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2171_5 ( .OUT(na2171_2), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2171_2_i) );
// C_AND/D///      x101y72     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2172_1 ( .OUT(na2172_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2172_2 ( .OUT(na2172_1), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2172_1_i) );
// C_///AND/D      x103y97     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2173_4 ( .OUT(na2173_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2173_5 ( .OUT(na2173_2), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2173_2_i) );
// C_AND/D///      x92y70     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2174_1 ( .OUT(na2174_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2174_2 ( .OUT(na2174_1), .CLK(1'b0), .EN(na1421_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2174_1_i) );
// C_///AND/D      x109y108     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2175_4 ( .OUT(na2175_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2175_5 ( .OUT(na2175_2), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2175_2_i) );
// C_AND/D///      x125y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2176_1 ( .OUT(na2176_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2176_2 ( .OUT(na2176_1), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2176_1_i) );
// C_///AND/D      x107y106     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2177_4 ( .OUT(na2177_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2177_5 ( .OUT(na2177_2), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2177_2_i) );
// C_AND/D///      x102y109     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2178_1 ( .OUT(na2178_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2178_2 ( .OUT(na2178_1), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2178_1_i) );
// C_///AND/D      x93y88     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2179_4 ( .OUT(na2179_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2179_5 ( .OUT(na2179_2), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2179_2_i) );
// C_AND/D///      x101y70     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2180_1 ( .OUT(na2180_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2180_2 ( .OUT(na2180_1), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2180_1_i) );
// C_///AND/D      x105y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2181_4 ( .OUT(na2181_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2181_5 ( .OUT(na2181_2), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2181_2_i) );
// C_AND/D///      x90y77     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2182_1 ( .OUT(na2182_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2182_2 ( .OUT(na2182_1), .CLK(1'b0), .EN(na1422_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2182_1_i) );
// C_///AND/D      x93y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2183_4 ( .OUT(na2183_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2183_5 ( .OUT(na2183_2), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2183_2_i) );
// C_AND/D///      x122y106     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2184_1 ( .OUT(na2184_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2184_2 ( .OUT(na2184_1), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2184_1_i) );
// C_///AND/D      x103y107     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2185_4 ( .OUT(na2185_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2185_5 ( .OUT(na2185_2), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2185_2_i) );
// C_AND/D///      x97y114     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2186_1 ( .OUT(na2186_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2186_2 ( .OUT(na2186_1), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2186_1_i) );
// C_///AND/D      x91y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2187_4 ( .OUT(na2187_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2187_5 ( .OUT(na2187_2), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2187_2_i) );
// C_AND/D///      x96y80     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2188_1 ( .OUT(na2188_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2188_2 ( .OUT(na2188_1), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2188_1_i) );
// C_///AND/D      x93y96     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2189_4 ( .OUT(na2189_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2189_5 ( .OUT(na2189_2), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2189_2_i) );
// C_AND/D///      x89y82     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2190_1 ( .OUT(na2190_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2190_2 ( .OUT(na2190_1), .CLK(1'b0), .EN(na1423_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2190_1_i) );
// C_///AND/D      x93y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2191_4 ( .OUT(na2191_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2191_5 ( .OUT(na2191_2), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2191_2_i) );
// C_AND/D///      x109y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2192_1 ( .OUT(na2192_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2192_2 ( .OUT(na2192_1), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2192_1_i) );
// C_///AND/D      x103y98     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2193_4 ( .OUT(na2193_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2193_5 ( .OUT(na2193_2), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2193_2_i) );
// C_AND/D///      x93y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2194_1 ( .OUT(na2194_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2194_2 ( .OUT(na2194_1), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2194_1_i) );
// C_///AND/D      x87y79     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2195_4 ( .OUT(na2195_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2195_5 ( .OUT(na2195_2), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2195_2_i) );
// C_AND/D///      x93y80     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2196_1 ( .OUT(na2196_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2196_2 ( .OUT(na2196_1), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2196_1_i) );
// C_///AND/D      x91y86     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2197_4 ( .OUT(na2197_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2197_5 ( .OUT(na2197_2), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2197_2_i) );
// C_AND/D///      x95y70     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2198_1 ( .OUT(na2198_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2198_2 ( .OUT(na2198_1), .CLK(1'b0), .EN(na1424_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2198_1_i) );
// C_///AND/D      x101y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2199_4 ( .OUT(na2199_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2199_5 ( .OUT(na2199_2), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2199_2_i) );
// C_AND/D///      x123y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2200_1 ( .OUT(na2200_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2200_2 ( .OUT(na2200_1), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2200_1_i) );
// C_///AND/D      x116y104     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2201_4 ( .OUT(na2201_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2201_5 ( .OUT(na2201_2), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2201_2_i) );
// C_AND/D///      x95y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2202_1 ( .OUT(na2202_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2202_2 ( .OUT(na2202_1), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2202_1_i) );
// C_///AND/D      x103y94     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2203_4 ( .OUT(na2203_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2203_5 ( .OUT(na2203_2), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2203_2_i) );
// C_AND/D///      x99y79     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2204_1 ( .OUT(na2204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2204_2 ( .OUT(na2204_1), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2204_1_i) );
// C_///AND/D      x101y92     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2205_4 ( .OUT(na2205_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2205_5 ( .OUT(na2205_2), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2205_2_i) );
// C_AND/D///      x87y70     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2206_1 ( .OUT(na2206_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2206_2 ( .OUT(na2206_1), .CLK(1'b0), .EN(na1425_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2206_1_i) );
// C_///AND/D      x107y112     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2207_4 ( .OUT(na2207_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2207_5 ( .OUT(na2207_2), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2207_2_i) );
// C_AND/D///      x124y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2208_1 ( .OUT(na2208_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2208_2 ( .OUT(na2208_1), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2208_1_i) );
// C_///AND/D      x109y110     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2209_4 ( .OUT(na2209_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2209_5 ( .OUT(na2209_2), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2209_2_i) );
// C_///AND/D      x105y114     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2210_4 ( .OUT(na2210_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2210_5 ( .OUT(na2210_2), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2210_2_i) );
// C_AND/D///      x104y92     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2211_1 ( .OUT(na2211_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2211_2 ( .OUT(na2211_1), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2211_1_i) );
// C_///AND/D      x95y67     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2212_4 ( .OUT(na2212_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2212_5 ( .OUT(na2212_2), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2212_2_i) );
// C_AND/D///      x102y87     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2213_1 ( .OUT(na2213_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2213_2 ( .OUT(na2213_1), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2213_1_i) );
// C_///AND/D      x93y74     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2214_4 ( .OUT(na2214_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2214_5 ( .OUT(na2214_2), .CLK(1'b0), .EN(na1426_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2214_2_i) );
// C_AND/D///      x91y108     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2215_1 ( .OUT(na2215_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2215_2 ( .OUT(na2215_1), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2215_1_i) );
// C_///AND/D      x119y107     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2216_4 ( .OUT(na2216_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2216_5 ( .OUT(na2216_2), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2216_2_i) );
// C_AND/D///      x104y96     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2217_1 ( .OUT(na2217_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2217_2 ( .OUT(na2217_1), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2217_1_i) );
// C_///AND/D      x91y111     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2218_4 ( .OUT(na2218_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2218_5 ( .OUT(na2218_2), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2218_2_i) );
// C_AND/D///      x93y94     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2219_1 ( .OUT(na2219_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2219_2 ( .OUT(na2219_1), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2219_1_i) );
// C_///AND/D      x93y70     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2220_4 ( .OUT(na2220_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2220_5 ( .OUT(na2220_2), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2220_2_i) );
// C_AND/D///      x99y90     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2221_1 ( .OUT(na2221_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2221_2 ( .OUT(na2221_1), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2221_1_i) );
// C_///AND/D      x91y66     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2222_4 ( .OUT(na2222_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2222_5 ( .OUT(na2222_2), .CLK(1'b0), .EN(na1427_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2222_2_i) );
// C_AND/D///      x105y110     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2223_1 ( .OUT(na2223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2223_2 ( .OUT(na2223_1), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2223_1_i) );
// C_AND/D///      x127y102     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2224_1 ( .OUT(na2224_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2224_2 ( .OUT(na2224_1), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2224_1_i) );
// C_AND/D///      x105y107     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2225_1 ( .OUT(na2225_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2225_2 ( .OUT(na2225_1), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2225_1_i) );
// C_///AND/D      x104y113     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2226_4 ( .OUT(na2226_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2226_5 ( .OUT(na2226_2), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2226_2_i) );
// C_AND/D///      x97y91     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2227_1 ( .OUT(na2227_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2227_2 ( .OUT(na2227_1), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2227_1_i) );
// C_///AND/D      x96y65     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2228_4 ( .OUT(na2228_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2228_5 ( .OUT(na2228_2), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2228_2_i) );
// C_AND/D///      x100y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2229_1 ( .OUT(na2229_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2229_2 ( .OUT(na2229_1), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2229_1_i) );
// C_///AND/D      x89y77     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2230_4 ( .OUT(na2230_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2230_5 ( .OUT(na2230_2), .CLK(1'b0), .EN(na1428_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2230_2_i) );
// C_AND/D///      x95y114     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2231_1 ( .OUT(na2231_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2231_2 ( .OUT(na2231_1), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2231_1_i) );
// C_///AND/D      x126y105     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2232_4 ( .OUT(na2232_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2232_5 ( .OUT(na2232_2), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2232_2_i) );
// C_AND/D///      x99y111     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2233_1 ( .OUT(na2233_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2233_2 ( .OUT(na2233_1), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2233_1_i) );
// C_///AND/D      x104y107     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2234_4 ( .OUT(na2234_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2234_5 ( .OUT(na2234_2), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2234_2_i) );
// C_AND/D///      x91y101     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2235_1 ( .OUT(na2235_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2235_2 ( .OUT(na2235_1), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2235_1_i) );
// C_///AND/D      x95y72     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2236_4 ( .OUT(na2236_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2236_5 ( .OUT(na2236_2), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2236_2_i) );
// C_AND/D///      x93y95     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2237_1 ( .OUT(na2237_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2237_2 ( .OUT(na2237_1), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2237_1_i) );
// C_///AND/D      x91y80     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2238_4 ( .OUT(na2238_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2238_5 ( .OUT(na2238_2), .CLK(1'b0), .EN(na1429_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2238_2_i) );
// C_AND/D///      x89y108     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2239_1 ( .OUT(na2239_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2239_2 ( .OUT(na2239_1), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2239_1_i) );
// C_///AND/D      x113y108     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2240_4 ( .OUT(na2240_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2240_5 ( .OUT(na2240_2), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2240_2_i) );
// C_AND/D///      x97y98     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2241_1 ( .OUT(na2241_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2241_2 ( .OUT(na2241_1), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2241_1_i) );
// C_///AND/D      x90y110     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2242_4 ( .OUT(na2242_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2242_5 ( .OUT(na2242_2), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2242_2_i) );
// C_AND/D///      x89y89     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2243_1 ( .OUT(na2243_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2243_2 ( .OUT(na2243_1), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2243_1_i) );
// C_///AND/D      x101y68     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2244_4 ( .OUT(na2244_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2244_5 ( .OUT(na2244_2), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2244_2_i) );
// C_AND/D///      x93y91     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2245_1 ( .OUT(na2245_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2245_2 ( .OUT(na2245_1), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2245_1_i) );
// C_///AND/D      x91y65     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2246_4 ( .OUT(na2246_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2246_5 ( .OUT(na2246_2), .CLK(1'b0), .EN(na1430_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2246_2_i) );
// C_AND/D///      x97y111     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2247_1 ( .OUT(na2247_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2247_2 ( .OUT(na2247_1), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2247_1_i) );
// C_///AND/D      x128y107     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2248_4 ( .OUT(na2248_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2248_5 ( .OUT(na2248_2), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2248_2_i) );
// C_AND/D///      x108y105     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2249_1 ( .OUT(na2249_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2249_2 ( .OUT(na2249_1), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2249_1_i) );
// C_///AND/D      x105y118     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2250_4 ( .OUT(na2250_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2250_5 ( .OUT(na2250_2), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2250_2_i) );
// C_AND/D///      x105y98     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2251_1 ( .OUT(na2251_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2251_2 ( .OUT(na2251_1), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2251_1_i) );
// C_///AND/D      x101y66     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2252_4 ( .OUT(na2252_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2252_5 ( .OUT(na2252_2), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2252_2_i) );
// C_///AND/D      x96y94     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2253_4 ( .OUT(na2253_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2253_5 ( .OUT(na2253_2), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2253_2_i) );
// C_///AND/D      x93y68     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2254_4 ( .OUT(na2254_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2254_5 ( .OUT(na2254_2), .CLK(1'b0), .EN(na1431_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2254_2_i) );
// C_AND/D///      x102y110     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2255_1 ( .OUT(na2255_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2255_2 ( .OUT(na2255_1), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2255_1_i) );
// C_///AND/D      x123y107     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2256_4 ( .OUT(na2256_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2256_5 ( .OUT(na2256_2), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2256_2_i) );
// C_AND/D///      x103y108     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2257_1 ( .OUT(na2257_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2257_2 ( .OUT(na2257_1), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2257_1_i) );
// C_///AND/D      x103y118     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2258_4 ( .OUT(na2258_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2258_5 ( .OUT(na2258_2), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2258_2_i) );
// C_AND/D///      x99y88     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2259_1 ( .OUT(na2259_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2259_2 ( .OUT(na2259_1), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2259_1_i) );
// C_///AND/D      x95y65     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2260_4 ( .OUT(na2260_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2260_5 ( .OUT(na2260_2), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2260_2_i) );
// C_AND/D///      x102y88     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2261_1 ( .OUT(na2261_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2261_2 ( .OUT(na2261_1), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2261_1_i) );
// C_///AND/D      x91y76     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2262_4 ( .OUT(na2262_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2262_5 ( .OUT(na2262_2), .CLK(1'b0), .EN(na1432_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2262_2_i) );
// C_AND/D///      x93y111     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2263_1 ( .OUT(na2263_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2263_2 ( .OUT(na2263_1), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2263_1_i) );
// C_///AND/D      x122y108     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2264_4 ( .OUT(na2264_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2264_5 ( .OUT(na2264_2), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2264_2_i) );
// C_AND/D///      x102y108     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2265_1 ( .OUT(na2265_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2265_2 ( .OUT(na2265_1), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2265_1_i) );
// C_///AND/D      x93y111     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2266_4 ( .OUT(na2266_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2266_5 ( .OUT(na2266_2), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2266_2_i) );
// C_AND/D///      x91y100     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2267_1 ( .OUT(na2267_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2267_2 ( .OUT(na2267_1), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2267_1_i) );
// C_///AND/D      x93y76     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2268_4 ( .OUT(na2268_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2268_5 ( .OUT(na2268_2), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2268_2_i) );
// C_AND/D///      x94y96     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2269_1 ( .OUT(na2269_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2269_2 ( .OUT(na2269_1), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2269_1_i) );
// C_///AND/D      x85y78     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2270_4 ( .OUT(na2270_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2270_5 ( .OUT(na2270_2), .CLK(1'b0), .EN(na1433_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2270_2_i) );
// C_AND/D///      x99y112     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2271_1 ( .OUT(na2271_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2271_2 ( .OUT(na2271_1), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2271_1_i) );
// C_///AND/D      x129y107     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2272_4 ( .OUT(na2272_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2272_5 ( .OUT(na2272_2), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2272_2_i) );
// C_AND/D///      x109y106     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2273_1 ( .OUT(na2273_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2273_2 ( .OUT(na2273_1), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2273_1_i) );
// C_///AND/D      x99y112     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2274_4 ( .OUT(na2274_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2274_5 ( .OUT(na2274_2), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2274_2_i) );
// C_AND/D///      x101y95     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2275_1 ( .OUT(na2275_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2275_2 ( .OUT(na2275_1), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2275_1_i) );
// C_///AND/D      x98y69     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2276_4 ( .OUT(na2276_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2276_5 ( .OUT(na2276_2), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2276_2_i) );
// C_AND/D///      x99y98     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2277_1 ( .OUT(na2277_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2277_2 ( .OUT(na2277_1), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2277_1_i) );
// C_///AND/D      x89y68     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2278_4 ( .OUT(na2278_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2278_5 ( .OUT(na2278_2), .CLK(1'b0), .EN(na1434_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2278_2_i) );
// C_AND/D///      x88y106     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2279_1 ( .OUT(na2279_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na735_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2279_2 ( .OUT(na2279_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2279_1_i) );
// C_///AND/D      x111y106     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2280_4 ( .OUT(na2280_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na736_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2280_5 ( .OUT(na2280_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2280_2_i) );
// C_AND/D///      x98y88     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2281_1 ( .OUT(na2281_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na737_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2281_2 ( .OUT(na2281_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2281_1_i) );
// C_///AND/D      x91y113     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2282_4 ( .OUT(na2282_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na738_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2282_5 ( .OUT(na2282_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2282_2_i) );
// C_///AND/D      x83y81     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2283_4 ( .OUT(na2283_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na739_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2283_5 ( .OUT(na2283_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2283_2_i) );
// C_///AND/D      x91y74     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2284_4 ( .OUT(na2284_2_i), .IN1(1'b1), .IN2(na740_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2284_5 ( .OUT(na2284_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2284_2_i) );
// C_AND/D///      x94y90     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2285_1 ( .OUT(na2285_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na741_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2285_2 ( .OUT(na2285_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2285_1_i) );
// C_///AND/D      x98y67     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2286_4 ( .OUT(na2286_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na742_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2286_5 ( .OUT(na2286_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2286_2_i) );
// C_AND/D///      x114y115     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2287_1 ( .OUT(na2287_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na743_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2287_2 ( .OUT(na2287_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2287_1_i) );
// C_///AND/D      x136y104     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2288_4 ( .OUT(na2288_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na744_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2288_5 ( .OUT(na2288_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2288_2_i) );
// C_AND/D///      x127y108     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2289_1 ( .OUT(na2289_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na745_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2289_2 ( .OUT(na2289_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2289_1_i) );
// C_///AND/D      x115y110     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2290_4 ( .OUT(na2290_2_i), .IN1(1'b1), .IN2(na746_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2290_5 ( .OUT(na2290_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2290_2_i) );
// C_AND/D///      x119y99     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2291_1 ( .OUT(na2291_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na747_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2291_2 ( .OUT(na2291_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2291_1_i) );
// C_///AND/D      x104y67     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2292_4 ( .OUT(na2292_2_i), .IN1(1'b1), .IN2(na748_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2292_5 ( .OUT(na2292_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2292_2_i) );
// C_AND/D///      x104y104     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2293_1 ( .OUT(na2293_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na749_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2293_2 ( .OUT(na2293_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2293_1_i) );
// C_///AND/D      x94y69     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2294_4 ( .OUT(na2294_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na750_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2294_5 ( .OUT(na2294_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2294_2_i) );
// C_AND/D///      x130y103     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2295_1 ( .OUT(na2295_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na751_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2295_2 ( .OUT(na2295_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2295_1_i) );
// C_///AND/D      x137y100     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2296_4 ( .OUT(na2296_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na752_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2296_5 ( .OUT(na2296_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2296_2_i) );
// C_AND/D///      x113y114     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2297_1 ( .OUT(na2297_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na753_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2297_2 ( .OUT(na2297_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2297_1_i) );
// C_///AND/D      x126y108     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2298_4 ( .OUT(na2298_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na754_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2298_5 ( .OUT(na2298_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2298_2_i) );
// C_AND/D///      x109y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2299_1 ( .OUT(na2299_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na755_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2299_2 ( .OUT(na2299_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2299_1_i) );
// C_///AND/D      x103y71     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2300_4 ( .OUT(na2300_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na756_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2300_5 ( .OUT(na2300_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2300_2_i) );
// C_AND/D///      x119y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2301_1 ( .OUT(na2301_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na757_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2301_2 ( .OUT(na2301_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2301_1_i) );
// C_///AND/D      x87y74     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2302_4 ( .OUT(na2302_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na758_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2302_5 ( .OUT(na2302_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2302_2_i) );
// C_AND/D///      x96y115     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2303_1 ( .OUT(na2303_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na759_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2303_2 ( .OUT(na2303_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2303_1_i) );
// C_///AND/D      x135y106     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2304_4 ( .OUT(na2304_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na760_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2304_5 ( .OUT(na2304_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2304_2_i) );
// C_AND/D///      x105y115     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2305_1 ( .OUT(na2305_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na761_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2305_2 ( .OUT(na2305_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2305_1_i) );
// C_///AND/D      x103y116     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2306_4 ( .OUT(na2306_2_i), .IN1(1'b1), .IN2(na762_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2306_5 ( .OUT(na2306_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2306_2_i) );
// C_AND/D///      x95y108     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2307_1 ( .OUT(na2307_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na763_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2307_2 ( .OUT(na2307_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2307_1_i) );
// C_///AND/D      x97y92     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2308_4 ( .OUT(na2308_2_i), .IN1(na764_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2308_5 ( .OUT(na2308_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2308_2_i) );
// C_AND/D///      x97y101     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2309_1 ( .OUT(na2309_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na765_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2309_2 ( .OUT(na2309_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2309_1_i) );
// C_///AND/D      x87y91     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2310_4 ( .OUT(na2310_2_i), .IN1(na766_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2310_5 ( .OUT(na2310_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2310_2_i) );
// C_AND/D///      x142y90     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2311_1 ( .OUT(na2311_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na807_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2311_2 ( .OUT(na2311_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2311_1_i) );
// C_AND/D///      x142y94     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2312_1 ( .OUT(na2312_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na852_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2312_2 ( .OUT(na2312_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2312_1_i) );
// C_AND/D///      x140y85     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2313_1 ( .OUT(na2313_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na862_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2313_2 ( .OUT(na2313_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2313_1_i) );
// C_///AND/D      x136y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2314_4 ( .OUT(na2314_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na866_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2314_5 ( .OUT(na2314_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2314_2_i) );
// C_AND/D///      x137y70     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2315_1 ( .OUT(na2315_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2315_2 ( .OUT(na2315_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2315_1_i) );
// C_///AND/D      x133y70     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2316_4 ( .OUT(na2316_2_i), .IN1(na875_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2316_5 ( .OUT(na2316_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2316_2_i) );
// C_AND/D///      x137y81     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2317_1 ( .OUT(na2317_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na877_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2317_2 ( .OUT(na2317_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2317_1_i) );
// C_///AND/D      x138y71     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2318_4 ( .OUT(na2318_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na881_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2318_5 ( .OUT(na2318_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2318_2_i) );
// C_AND/D///      x118y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2319_1 ( .OUT(na2319_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na215_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2319_2 ( .OUT(na2319_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2319_1_i) );
// C_///AND/D      x124y98     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2320_4 ( .OUT(na2320_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na263_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2320_5 ( .OUT(na2320_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2320_2_i) );
// C_AND/D///      x113y80     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2321_1 ( .OUT(na2321_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na275_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2321_2 ( .OUT(na2321_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2321_1_i) );
// C_///AND/D      x118y98     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2322_4 ( .OUT(na2322_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na281_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2322_5 ( .OUT(na2322_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2322_2_i) );
// C_AND/D///      x110y77     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2323_1 ( .OUT(na2323_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na293_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2323_2 ( .OUT(na2323_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2323_1_i) );
// C_///AND/D      x112y79     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2324_4 ( .OUT(na2324_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na298_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2324_5 ( .OUT(na2324_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2324_2_i) );
// C_AND/D///      x109y86     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2325_1 ( .OUT(na2325_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na308_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2325_2 ( .OUT(na2325_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2325_1_i) );
// C_///AND/D      x111y80     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2326_4 ( .OUT(na2326_2_i), .IN1(na312_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2326_5 ( .OUT(na2326_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2326_2_i) );
// C_AND/D///      x129y102     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2327_1 ( .OUT(na2327_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na959_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2327_2 ( .OUT(na2327_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2327_1_i) );
// C_///AND/D      x135y102     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2328_4 ( .OUT(na2328_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1003_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2328_5 ( .OUT(na2328_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2328_2_i) );
// C_AND/D///      x132y93     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2329_1 ( .OUT(na2329_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1012_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2329_2 ( .OUT(na2329_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2329_1_i) );
// C_///AND/D      x131y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2330_4 ( .OUT(na2330_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1019_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2330_5 ( .OUT(na2330_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2330_2_i) );
// C_AND/D///      x127y83     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2331_1 ( .OUT(na2331_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1025_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2331_2 ( .OUT(na2331_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2331_1_i) );
// C_///AND/D      x121y78     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2332_4 ( .OUT(na2332_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1029_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2332_5 ( .OUT(na2332_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2332_2_i) );
// C_AND/D///      x117y94     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2333_1 ( .OUT(na2333_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2333_2 ( .OUT(na2333_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2333_1_i) );
// C_///AND/D      x123y90     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2334_4 ( .OUT(na2334_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1034_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2334_5 ( .OUT(na2334_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2334_2_i) );
// C_AND/D///      x137y95     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2335_1 ( .OUT(na2335_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na884_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2335_2 ( .OUT(na2335_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2335_1_i) );
// C_///AND/D      x138y96     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2336_4 ( .OUT(na2336_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na926_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2336_5 ( .OUT(na2336_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2336_2_i) );
// C_AND/D///      x134y82     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2337_1 ( .OUT(na2337_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na935_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2337_2 ( .OUT(na2337_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2337_1_i) );
// C_///AND/D      x138y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2338_4 ( .OUT(na2338_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na941_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2338_5 ( .OUT(na2338_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2338_2_i) );
// C_AND/D///      x129y70     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2339_1 ( .OUT(na2339_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2339_2 ( .OUT(na2339_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2339_1_i) );
// C_///AND/D      x129y70     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2340_4 ( .OUT(na2340_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na952_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2340_5 ( .OUT(na2340_2), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2340_2_i) );
// C_AND/D///      x133y78     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2341_1 ( .OUT(na2341_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na955_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2341_2 ( .OUT(na2341_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2341_1_i) );
// C_AND/D///      x131y70     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2342_1 ( .OUT(na2342_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na957_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2342_2 ( .OUT(na2342_1), .CLK(1'b0), .EN(na323_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2342_1_i) );
// C_AND/D///      x141y94     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2343_1 ( .OUT(na2343_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na884_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2343_2 ( .OUT(na2343_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2343_1_i) );
// C_///AND/D      x141y95     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2344_4 ( .OUT(na2344_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na926_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2344_5 ( .OUT(na2344_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2344_2_i) );
// C_AND/D///      x140y73     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2345_1 ( .OUT(na2345_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na935_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2345_2 ( .OUT(na2345_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2345_1_i) );
// C_///AND/D      x142y92     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2346_4 ( .OUT(na2346_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na941_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2346_5 ( .OUT(na2346_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2346_2_i) );
// C_AND/D///      x137y66     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2347_1 ( .OUT(na2347_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2347_2 ( .OUT(na2347_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2347_1_i) );
// C_///AND/D      x136y67     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2348_4 ( .OUT(na2348_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na952_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2348_5 ( .OUT(na2348_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2348_2_i) );
// C_AND/D///      x139y72     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2349_1 ( .OUT(na2349_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na955_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2349_2 ( .OUT(na2349_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2349_1_i) );
// C_///AND/D      x137y65     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2350_4 ( .OUT(na2350_2_i), .IN1(na957_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2350_5 ( .OUT(na2350_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2350_2_i) );
// C_AND/D///      x139y94     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2351_1 ( .OUT(na2351_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na807_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2351_2 ( .OUT(na2351_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2351_1_i) );
// C_///AND/D      x144y102     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2352_4 ( .OUT(na2352_2_i), .IN1(na852_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2352_5 ( .OUT(na2352_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2352_2_i) );
// C_AND/D///      x141y88     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2353_1 ( .OUT(na2353_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na862_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2353_2 ( .OUT(na2353_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2353_1_i) );
// C_///AND/D      x134y91     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2354_4 ( .OUT(na2354_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na866_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2354_5 ( .OUT(na2354_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2354_2_i) );
// C_AND/D///      x140y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2355_1 ( .OUT(na2355_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2355_2 ( .OUT(na2355_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2355_1_i) );
// C_///AND/D      x127y72     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2356_4 ( .OUT(na2356_2_i), .IN1(na875_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2356_5 ( .OUT(na2356_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2356_2_i) );
// C_AND/D///      x135y86     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2357_1 ( .OUT(na2357_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na877_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2357_2 ( .OUT(na2357_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2357_1_i) );
// C_///AND/D      x129y74     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2358_4 ( .OUT(na2358_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na881_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2358_5 ( .OUT(na2358_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2358_2_i) );
// C_AND/D///      x118y92     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2359_1 ( .OUT(na2359_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na215_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2359_2 ( .OUT(na2359_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2359_1_i) );
// C_///AND/D      x113y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2360_4 ( .OUT(na2360_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na263_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2360_5 ( .OUT(na2360_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2360_2_i) );
// C_AND/D///      x114y83     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2361_1 ( .OUT(na2361_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na275_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2361_2 ( .OUT(na2361_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2361_1_i) );
// C_///AND/D      x115y102     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2362_4 ( .OUT(na2362_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na281_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2362_5 ( .OUT(na2362_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2362_2_i) );
// C_AND/D///      x115y81     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2363_1 ( .OUT(na2363_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na293_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2363_2 ( .OUT(na2363_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2363_1_i) );
// C_///AND/D      x118y84     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2364_4 ( .OUT(na2364_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na298_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2364_5 ( .OUT(na2364_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2364_2_i) );
// C_AND/D///      x112y89     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2365_1 ( .OUT(na2365_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na308_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2365_2 ( .OUT(na2365_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2365_1_i) );
// C_///AND/D      x111y76     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2366_4 ( .OUT(na2366_2_i), .IN1(na312_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2366_5 ( .OUT(na2366_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2366_2_i) );
// C_AND/D///      x131y102     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2367_1 ( .OUT(na2367_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na959_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2367_2 ( .OUT(na2367_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2367_1_i) );
// C_///AND/D      x133y101     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2368_4 ( .OUT(na2368_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1003_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2368_5 ( .OUT(na2368_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2368_2_i) );
// C_AND/D///      x127y92     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2369_1 ( .OUT(na2369_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1012_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2369_2 ( .OUT(na2369_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2369_1_i) );
// C_///AND/D      x134y93     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2370_4 ( .OUT(na2370_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1019_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2370_5 ( .OUT(na2370_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2370_2_i) );
// C_///AND/D      x131y90     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2371_4 ( .OUT(na2371_2_i), .IN1(na1025_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2371_5 ( .OUT(na2371_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2371_2_i) );
// C_///AND/D      x122y77     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2372_4 ( .OUT(na2372_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1029_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2372_5 ( .OUT(na2372_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2372_2_i) );
// C_AND/D///      x120y95     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2373_1 ( .OUT(na2373_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2373_2 ( .OUT(na2373_1), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2373_1_i) );
// C_///AND/D      x128y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2374_4 ( .OUT(na2374_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1034_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2374_5 ( .OUT(na2374_2), .CLK(1'b0), .EN(na27_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2374_2_i) );
// C_AND/D///      x135y98     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2375_1 ( .OUT(na2375_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na959_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2375_2 ( .OUT(na2375_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2375_1_i) );
// C_///AND/D      x140y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2376_4 ( .OUT(na2376_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1003_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2376_5 ( .OUT(na2376_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2376_2_i) );
// C_AND/D///      x133y90     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2377_1 ( .OUT(na2377_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1012_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2377_2 ( .OUT(na2377_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2377_1_i) );
// C_///AND/D      x131y96     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2378_4 ( .OUT(na2378_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1019_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2378_5 ( .OUT(na2378_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2378_2_i) );
// C_AND/D///      x141y76     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2379_1 ( .OUT(na2379_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1025_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2379_2 ( .OUT(na2379_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2379_1_i) );
// C_///AND/D      x129y73     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2380_4 ( .OUT(na2380_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1029_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2380_5 ( .OUT(na2380_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2380_2_i) );
// C_AND/D///      x125y91     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2381_1 ( .OUT(na2381_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2381_2 ( .OUT(na2381_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2381_1_i) );
// C_///AND/D      x129y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2382_4 ( .OUT(na2382_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1034_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2382_5 ( .OUT(na2382_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2382_2_i) );
// C_AND/D///      x140y97     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2383_1 ( .OUT(na2383_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na884_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2383_2 ( .OUT(na2383_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2383_1_i) );
// C_///AND/D      x140y95     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2384_4 ( .OUT(na2384_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na926_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2384_5 ( .OUT(na2384_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2384_2_i) );
// C_AND/D///      x139y80     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2385_1 ( .OUT(na2385_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na935_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2385_2 ( .OUT(na2385_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2385_1_i) );
// C_///AND/D      x145y88     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2386_4 ( .OUT(na2386_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na941_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2386_5 ( .OUT(na2386_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2386_2_i) );
// C_AND/D///      x135y68     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2387_1 ( .OUT(na2387_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2387_2 ( .OUT(na2387_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2387_1_i) );
// C_///AND/D      x129y68     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2388_4 ( .OUT(na2388_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na952_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2388_5 ( .OUT(na2388_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2388_2_i) );
// C_AND/D///      x136y73     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2389_1 ( .OUT(na2389_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na955_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2389_2 ( .OUT(na2389_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2389_1_i) );
// C_///AND/D      x136y68     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2390_4 ( .OUT(na2390_2_i), .IN1(na957_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2390_5 ( .OUT(na2390_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2390_2_i) );
// C_AND/D///      x135y94     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2391_1 ( .OUT(na2391_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na807_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2391_2 ( .OUT(na2391_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2391_1_i) );
// C_///AND/D      x138y101     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2392_4 ( .OUT(na2392_2_i), .IN1(na852_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2392_5 ( .OUT(na2392_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2392_2_i) );
// C_AND/D///      x136y89     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2393_1 ( .OUT(na2393_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na862_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2393_2 ( .OUT(na2393_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2393_1_i) );
// C_///AND/D      x133y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2394_4 ( .OUT(na2394_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na866_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2394_5 ( .OUT(na2394_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2394_2_i) );
// C_AND/D///      x136y79     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2395_1 ( .OUT(na2395_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2395_2 ( .OUT(na2395_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2395_1_i) );
// C_///AND/D      x127y75     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2396_4 ( .OUT(na2396_2_i), .IN1(na875_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2396_5 ( .OUT(na2396_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2396_2_i) );
// C_AND/D///      x134y88     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2397_1 ( .OUT(na2397_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na877_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2397_2 ( .OUT(na2397_1), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2397_1_i) );
// C_///AND/D      x131y82     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2398_4 ( .OUT(na2398_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na881_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2398_5 ( .OUT(na2398_2), .CLK(1'b0), .EN(na1437_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2398_2_i) );
// C_AND/D///      x150y74     80'h40_F800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2399_1 ( .OUT(na2399_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1349_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2399_2 ( .OUT(na2399_1), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2399_1_i) );
// C_///AND/D      x149y89     80'h40_F800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2400_4 ( .OUT(na2400_2_i), .IN1(na1350_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2400_5 ( .OUT(na2400_2), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2400_2_i) );
// C_///AND/D      x146y89     80'h40_F800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2401_4 ( .OUT(na2401_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1351_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2401_5 ( .OUT(na2401_2), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2401_2_i) );
// C_///AND/D      x149y95     80'h40_F800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2402_4 ( .OUT(na2402_2_i), .IN1(1'b1), .IN2(na1352_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2402_5 ( .OUT(na2402_2), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2402_2_i) );
// C_AND/D///      x148y92     80'h40_F800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2403_1 ( .OUT(na2403_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1353_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2403_2 ( .OUT(na2403_1), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2403_1_i) );
// C_///AND/D      x148y92     80'h40_F800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2404_4 ( .OUT(na2404_2_i), .IN1(1'b1), .IN2(na1354_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2404_5 ( .OUT(na2404_2), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2404_2_i) );
// C_AND/D///      x147y92     80'h40_F800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2405_1 ( .OUT(na2405_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1355_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2405_2 ( .OUT(na2405_1), .CLK(1'b0), .EN(na1382_2), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2405_1_i) );
// C_///AND/D      x138y76     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2406_4 ( .OUT(na2406_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1125_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2406_5 ( .OUT(na2406_2), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2406_2_i) );
// C_AND/D///      x135y84     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2407_1 ( .OUT(na2407_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1127_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2407_2 ( .OUT(na2407_1), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2407_1_i) );
// C_///AND/D      x136y70     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2408_4 ( .OUT(na2408_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1128_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2408_5 ( .OUT(na2408_2), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2408_2_i) );
// C_AND/D///      x132y85     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2409_1 ( .OUT(na2409_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1129_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2409_2 ( .OUT(na2409_1), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2409_1_i) );
// C_///AND/D      x133y71     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2410_4 ( .OUT(na2410_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1130_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2410_5 ( .OUT(na2410_2), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2410_2_i) );
// C_AND/D///      x133y71     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2411_1 ( .OUT(na2411_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1131_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2411_2 ( .OUT(na2411_1), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2411_1_i) );
// C_///AND/D      x136y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2412_4 ( .OUT(na2412_2_i), .IN1(1'b1), .IN2(na1132_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2412_5 ( .OUT(na2412_2), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2412_2_i) );
// C_AND/D///      x132y70     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2413_1 ( .OUT(na2413_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1133_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2413_2 ( .OUT(na2413_1), .CLK(1'b0), .EN(na322_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2413_1_i) );
// C_///AND/D      x125y73     80'h40_E400_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2415_4 ( .OUT(na2415_2_i), .IN1(1'b1), .IN2(na1320_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2415_5 ( .OUT(na2415_2), .CLK(1'b0), .EN(~na21_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2415_2_i) );
// C_AND/D//AND/D      x115y90     80'h40_E400_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2416_1 ( .OUT(na2416_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1321_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2416_2 ( .OUT(na2416_1), .CLK(1'b0), .EN(~na21_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2416_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2416_4 ( .OUT(na2416_2_i), .IN1(na1319_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2416_5 ( .OUT(na2416_2), .CLK(1'b0), .EN(~na21_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2416_2_i) );
// C_AND/D///      x122y71     80'h40_E400_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2417_1 ( .OUT(na2417_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1322_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2417_2 ( .OUT(na2417_1), .CLK(1'b0), .EN(~na21_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2417_1_i) );
// C_///AND/D      x96y103     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2418_4 ( .OUT(na2418_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na542_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2418_5 ( .OUT(na2418_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2418_2_i) );
// C_AND/D///      x110y99     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2419_1 ( .OUT(na2419_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na544_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2419_2 ( .OUT(na2419_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2419_1_i) );
// C_///AND/D      x107y81     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2420_4 ( .OUT(na2420_2_i), .IN1(na545_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2420_5 ( .OUT(na2420_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2420_2_i) );
// C_AND/D///      x95y107     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2421_1 ( .OUT(na2421_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na546_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2421_2 ( .OUT(na2421_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2421_1_i) );
// C_///AND/D      x91y78     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2422_4 ( .OUT(na2422_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na547_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2422_5 ( .OUT(na2422_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2422_2_i) );
// C_AND/D///      x103y86     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2423_1 ( .OUT(na2423_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2423_2 ( .OUT(na2423_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2423_1_i) );
// C_AND/D//AND/D      x96y88     80'h40_E800_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2424_1 ( .OUT(na2424_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na549_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2424_2 ( .OUT(na2424_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2424_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2424_4 ( .OUT(na2424_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na613_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2424_5 ( .OUT(na2424_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2424_2_i) );
// C_///AND/D      x103y69     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2425_4 ( .OUT(na2425_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na550_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2425_5 ( .OUT(na2425_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2425_2_i) );
// C_AND/D///      x112y109     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2426_1 ( .OUT(na2426_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na551_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2426_2 ( .OUT(na2426_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2426_1_i) );
// C_AND/D//AND/D      x132y101     80'h40_E800_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2427_1 ( .OUT(na2427_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na552_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2427_2 ( .OUT(na2427_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2427_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2427_4 ( .OUT(na2427_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na616_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2427_5 ( .OUT(na2427_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2427_2_i) );
// C_///AND/D      x122y100     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2428_4 ( .OUT(na2428_2_i), .IN1(1'b1), .IN2(na553_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2428_5 ( .OUT(na2428_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2428_2_i) );
// C_AND/D///      x110y108     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2429_1 ( .OUT(na2429_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na554_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2429_2 ( .OUT(na2429_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2429_1_i) );
// C_///AND/D      x120y93     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2430_4 ( .OUT(na2430_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na555_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2430_5 ( .OUT(na2430_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2430_2_i) );
// C_AND/D//AND/D      x110y76     80'h40_E800_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2431_1 ( .OUT(na2431_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na556_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2431_2 ( .OUT(na2431_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2431_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2431_4 ( .OUT(na2431_2_i), .IN1(1'b1), .IN2(na620_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2431_5 ( .OUT(na2431_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2431_2_i) );
// C_AND/D///      x109y97     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2432_1 ( .OUT(na2432_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na557_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2432_2 ( .OUT(na2432_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2432_1_i) );
// C_///AND/D      x102y73     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2433_4 ( .OUT(na2433_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na558_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2433_5 ( .OUT(na2433_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2433_2_i) );
// C_AND/D//AND/D      x129y104     80'h40_E800_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2434_1 ( .OUT(na2434_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na559_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2434_2 ( .OUT(na2434_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2434_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2434_4 ( .OUT(na2434_2_i), .IN1(1'b1), .IN2(na623_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2434_5 ( .OUT(na2434_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2434_2_i) );
// C_AND/D//AND/D      x133y99     80'h40_E800_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2435_1 ( .OUT(na2435_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na560_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2435_2 ( .OUT(na2435_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2435_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2435_4 ( .OUT(na2435_2_i), .IN1(na624_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2435_5 ( .OUT(na2435_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2435_2_i) );
// C_AND/D///      x118y106     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2436_1 ( .OUT(na2436_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na561_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2436_2 ( .OUT(na2436_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2436_1_i) );
// C_AND/D///      x117y109     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2437_1 ( .OUT(na2437_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na562_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2437_2 ( .OUT(na2437_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2437_1_i) );
// C_AND/D///      x116y92     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2438_1 ( .OUT(na2438_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na563_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2438_2 ( .OUT(na2438_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2438_1_i) );
// C_///AND/D      x105y65     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2439_4 ( .OUT(na2439_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na564_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2439_5 ( .OUT(na2439_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2439_2_i) );
// C_AND/D//AND/D      x116y83     80'h40_E800_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2440_1 ( .OUT(na2440_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na565_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2440_2 ( .OUT(na2440_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2440_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2440_4 ( .OUT(na2440_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na629_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2440_5 ( .OUT(na2440_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2440_2_i) );
// C_AND/D///      x102y83     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2441_1 ( .OUT(na2441_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na566_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2441_2 ( .OUT(na2441_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2441_1_i) );
// C_///AND/D      x111y104     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2442_4 ( .OUT(na2442_2_i), .IN1(na567_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2442_5 ( .OUT(na2442_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2442_2_i) );
// C_AND/D///      x127y103     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2443_1 ( .OUT(na2443_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na568_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2443_2 ( .OUT(na2443_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2443_1_i) );
// C_///AND/D      x117y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2444_4 ( .OUT(na2444_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na569_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2444_5 ( .OUT(na2444_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2444_2_i) );
// C_AND/D///      x105y109     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2445_1 ( .OUT(na2445_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na570_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2445_2 ( .OUT(na2445_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2445_1_i) );
// C_///AND/D      x101y104     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2446_4 ( .OUT(na2446_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na571_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2446_5 ( .OUT(na2446_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2446_2_i) );
// C_AND/D///      x102y90     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2447_1 ( .OUT(na2447_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na572_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2447_2 ( .OUT(na2447_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2447_1_i) );
// C_///AND/D      x100y95     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2448_4 ( .OUT(na2448_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na573_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2448_5 ( .OUT(na2448_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2448_2_i) );
// C_AND/D///      x102y93     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2449_1 ( .OUT(na2449_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na574_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2449_2 ( .OUT(na2449_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2449_1_i) );
// C_///AND/D      x99y107     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2450_4 ( .OUT(na2450_2_i), .IN1(1'b1), .IN2(na575_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2450_5 ( .OUT(na2450_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2450_2_i) );
// C_AND/D//AND/D      x130y105     80'h40_E800_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2451_1 ( .OUT(na2451_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na576_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2451_2 ( .OUT(na2451_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2451_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2451_4 ( .OUT(na2451_2_i), .IN1(na728_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2451_5 ( .OUT(na2451_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2451_2_i) );
// C_AND/D///      x110y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2452_1 ( .OUT(na2452_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na577_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2452_2 ( .OUT(na2452_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2452_1_i) );
// C_///AND/D      x116y112     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2453_4 ( .OUT(na2453_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na578_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2453_5 ( .OUT(na2453_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2453_2_i) );
// C_AND/D///      x100y98     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2454_1 ( .OUT(na2454_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na579_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2454_2 ( .OUT(na2454_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2454_1_i) );
// C_///AND/D      x100y83     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2455_4 ( .OUT(na2455_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na580_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2455_5 ( .OUT(na2455_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2455_2_i) );
// C_AND/D//AND/D      x95y100     80'h40_E800_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2456_1 ( .OUT(na2456_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na581_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2456_2 ( .OUT(na2456_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2456_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2456_4 ( .OUT(na2456_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na733_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2456_5 ( .OUT(na2456_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2456_2_i) );
// C_AND/D///      x101y90     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2457_1 ( .OUT(na2457_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na582_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2457_2 ( .OUT(na2457_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2457_1_i) );
// C_///AND/D      x97y105     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2458_4 ( .OUT(na2458_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na583_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2458_5 ( .OUT(na2458_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2458_2_i) );
// C_AND/D///      x115y105     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2459_1 ( .OUT(na2459_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na584_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2459_2 ( .OUT(na2459_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2459_1_i) );
// C_///AND/D      x108y81     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2460_4 ( .OUT(na2460_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na585_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2460_5 ( .OUT(na2460_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2460_2_i) );
// C_AND/D///      x98y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2461_1 ( .OUT(na2461_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na586_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2461_2 ( .OUT(na2461_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2461_1_i) );
// C_///AND/D      x97y81     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2462_4 ( .OUT(na2462_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2462_5 ( .OUT(na2462_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2462_2_i) );
// C_AND/D///      x105y79     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2463_1 ( .OUT(na2463_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na588_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2463_2 ( .OUT(na2463_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2463_1_i) );
// C_AND/D//AND/D      x99y92     80'h40_E800_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2464_1 ( .OUT(na2464_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na589_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2464_2 ( .OUT(na2464_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2464_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2464_4 ( .OUT(na2464_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na709_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2464_5 ( .OUT(na2464_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2464_2_i) );
// C_///AND/D      x102y67     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2465_4 ( .OUT(na2465_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na590_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2465_5 ( .OUT(na2465_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2465_2_i) );
// C_AND/D///      x116y112     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2466_1 ( .OUT(na2466_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na591_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2466_2 ( .OUT(na2466_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2466_1_i) );
// C_AND/D//AND/D      x135y104     80'h40_E800_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2467_1 ( .OUT(na2467_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na592_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2467_2 ( .OUT(na2467_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2467_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2467_4 ( .OUT(na2467_2_i), .IN1(1'b1), .IN2(na712_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2467_5 ( .OUT(na2467_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2467_2_i) );
// C_///AND/D      x121y99     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2468_4 ( .OUT(na2468_2_i), .IN1(na593_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2468_5 ( .OUT(na2468_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2468_2_i) );
// C_AND/D///      x111y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2469_1 ( .OUT(na2469_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na594_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2469_2 ( .OUT(na2469_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2469_1_i) );
// C_///AND/D      x120y96     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2470_4 ( .OUT(na2470_2_i), .IN1(1'b1), .IN2(na595_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2470_5 ( .OUT(na2470_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2470_2_i) );
// C_AND/D//AND/D      x107y72     80'h40_E800_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2471_1 ( .OUT(na2471_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na596_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2471_2 ( .OUT(na2471_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2471_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2471_4 ( .OUT(na2471_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na716_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2471_5 ( .OUT(na2471_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2471_2_i) );
// C_AND/D///      x112y95     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2472_1 ( .OUT(na2472_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na597_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2472_2 ( .OUT(na2472_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2472_1_i) );
// C_AND/D///      x107y71     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2473_1 ( .OUT(na2473_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na598_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2473_2 ( .OUT(na2473_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2473_1_i) );
// C_AND/D//AND/D      x125y103     80'h40_E800_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2474_1 ( .OUT(na2474_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na599_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2474_2 ( .OUT(na2474_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2474_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2474_4 ( .OUT(na2474_2_i), .IN1(1'b1), .IN2(na719_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2474_5 ( .OUT(na2474_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2474_2_i) );
// C_AND/D//AND/D      x136y99     80'h40_E800_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2475_1 ( .OUT(na2475_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na600_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2475_2 ( .OUT(na2475_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2475_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2475_4 ( .OUT(na2475_2_i), .IN1(1'b1), .IN2(na720_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2475_5 ( .OUT(na2475_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2475_2_i) );
// C_AND/D///      x116y107     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2476_1 ( .OUT(na2476_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na601_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2476_2 ( .OUT(na2476_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2476_1_i) );
// C_///AND/D      x122y109     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2477_4 ( .OUT(na2477_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na602_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2477_5 ( .OUT(na2477_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2477_2_i) );
// C_AND/D///      x111y91     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2478_1 ( .OUT(na2478_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na603_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2478_2 ( .OUT(na2478_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2478_1_i) );
// C_///AND/D      x107y74     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2479_4 ( .OUT(na2479_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na604_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2479_5 ( .OUT(na2479_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2479_2_i) );
// C_AND/D//AND/D      x117y87     80'h40_E800_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2480_1 ( .OUT(na2480_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na605_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2480_2 ( .OUT(na2480_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2480_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2480_4 ( .OUT(na2480_2_i), .IN1(1'b1), .IN2(na725_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2480_5 ( .OUT(na2480_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2480_2_i) );
// C_AND/D///      x99y83     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2481_1 ( .OUT(na2481_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na606_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2481_2 ( .OUT(na2481_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2481_1_i) );
// C_///AND/D      x88y101     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2482_4 ( .OUT(na2482_2_i), .IN1(na1480_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2482_5 ( .OUT(na2482_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2482_2_i) );
// C_AND/D///      x101y102     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2483_1 ( .OUT(na2483_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1481_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2483_2 ( .OUT(na2483_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2483_1_i) );
// C_///AND/D      x98y73     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2484_4 ( .OUT(na2484_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1482_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2484_5 ( .OUT(na2484_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2484_2_i) );
// C_AND/D///      x91y116     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2485_1 ( .OUT(na2485_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1483_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2485_2 ( .OUT(na2485_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2485_1_i) );
// C_///AND/D      x90y79     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2486_4 ( .OUT(na2486_2_i), .IN1(na1484_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2486_5 ( .OUT(na2486_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2486_2_i) );
// C_AND/D///      x93y85     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2487_1 ( .OUT(na2487_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1485_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2487_2 ( .OUT(na2487_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2487_1_i) );
// C_///AND/D      x88y86     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2488_4 ( .OUT(na2488_2_i), .IN1(1'b1), .IN2(na1486_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2488_5 ( .OUT(na2488_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2488_2_i) );
// C_AND/D///      x99y72     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2489_1 ( .OUT(na2489_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1487_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2489_2 ( .OUT(na2489_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2489_1_i) );
// C_///AND/D      x118y115     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2490_4 ( .OUT(na2490_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1488_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2490_5 ( .OUT(na2490_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2490_2_i) );
// C_AND/D///      x136y103     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2491_1 ( .OUT(na2491_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1489_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2491_2 ( .OUT(na2491_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2491_1_i) );
// C_///AND/D      x136y106     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2492_4 ( .OUT(na2492_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1490_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2492_5 ( .OUT(na2492_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2492_2_i) );
// C_AND/D///      x111y109     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2493_1 ( .OUT(na2493_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1491_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2493_2 ( .OUT(na2493_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2493_1_i) );
// C_///AND/D      x132y90     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2494_4 ( .OUT(na2494_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1492_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2494_5 ( .OUT(na2494_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2494_2_i) );
// C_AND/D///      x106y75     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2495_1 ( .OUT(na2495_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1493_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2495_2 ( .OUT(na2495_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2495_1_i) );
// C_///AND/D      x118y108     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2496_4 ( .OUT(na2496_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1494_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2496_5 ( .OUT(na2496_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2496_2_i) );
// C_AND/D///      x92y79     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2497_1 ( .OUT(na2497_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1495_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2497_2 ( .OUT(na2497_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2497_1_i) );
// C_///AND/D      x134y104     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2498_4 ( .OUT(na2498_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1496_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2498_5 ( .OUT(na2498_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2498_2_i) );
// C_AND/D///      x134y100     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2499_1 ( .OUT(na2499_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1497_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2499_2 ( .OUT(na2499_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2499_1_i) );
// C_///AND/D      x115y106     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2500_4 ( .OUT(na2500_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1498_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2500_5 ( .OUT(na2500_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2500_2_i) );
// C_AND/D///      x122y107     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2501_1 ( .OUT(na2501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1499_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2501_2 ( .OUT(na2501_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2501_1_i) );
// C_///AND/D      x111y78     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2502_4 ( .OUT(na2502_2_i), .IN1(1'b1), .IN2(na1500_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2502_5 ( .OUT(na2502_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2502_2_i) );
// C_AND/D///      x108y65     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2503_1 ( .OUT(na2503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1501_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2503_2 ( .OUT(na2503_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2503_1_i) );
// C_///AND/D      x117y78     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2504_4 ( .OUT(na2504_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1502_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2504_5 ( .OUT(na2504_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2504_2_i) );
// C_///AND/D      x96y79     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2505_4 ( .OUT(na2505_2_i), .IN1(1'b1), .IN2(na1503_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2505_5 ( .OUT(na2505_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2505_2_i) );
// C_///AND/D      x95y116     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2506_4 ( .OUT(na2506_2_i), .IN1(na1469_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2506_5 ( .OUT(na2506_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2506_2_i) );
// C_AND/D///      x124y108     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2507_1 ( .OUT(na2507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1470_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2507_2 ( .OUT(na2507_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2507_1_i) );
// C_///AND/D      x111y116     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2508_4 ( .OUT(na2508_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1471_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2508_5 ( .OUT(na2508_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2508_2_i) );
// C_AND/D///      x104y115     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2509_1 ( .OUT(na2509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1473_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2509_2 ( .OUT(na2509_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2509_1_i) );
// C_///AND/D      x107y109     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2510_4 ( .OUT(na2510_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1475_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2510_5 ( .OUT(na2510_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2510_2_i) );
// C_AND/D///      x89y101     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2511_1 ( .OUT(na2511_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1476_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2511_2 ( .OUT(na2511_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2511_1_i) );
// C_///AND/D      x103y111     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2512_4 ( .OUT(na2512_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1477_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2512_5 ( .OUT(na2512_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2512_2_i) );
// C_AND/D///      x96y106     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2513_1 ( .OUT(na2513_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1478_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2513_2 ( .OUT(na2513_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2513_1_i) );
// C_///AND/D      x91y110     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2514_4 ( .OUT(na2514_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1504_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2514_5 ( .OUT(na2514_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2514_2_i) );
// C_AND/D///      x100y107     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2515_1 ( .OUT(na2515_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1505_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2515_2 ( .OUT(na2515_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2515_1_i) );
// C_///AND/D      x91y73     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2516_4 ( .OUT(na2516_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1506_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2516_5 ( .OUT(na2516_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2516_2_i) );
// C_AND/D///      x89y115     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2517_1 ( .OUT(na2517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1507_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2517_2 ( .OUT(na2517_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2517_1_i) );
// C_///AND/D      x88y80     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2518_4 ( .OUT(na2518_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1508_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2518_5 ( .OUT(na2518_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2518_2_i) );
// C_AND/D///      x89y85     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2519_1 ( .OUT(na2519_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1509_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2519_2 ( .OUT(na2519_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2519_1_i) );
// C_///AND/D      x87y86     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2520_4 ( .OUT(na2520_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1510_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2520_5 ( .OUT(na2520_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2520_2_i) );
// C_AND/D///      x93y72     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2521_1 ( .OUT(na2521_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1511_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2521_2 ( .OUT(na2521_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2521_1_i) );
// C_///AND/D      x115y115     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2522_4 ( .OUT(na2522_2_i), .IN1(1'b1), .IN2(na1512_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2522_5 ( .OUT(na2522_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2522_2_i) );
// C_AND/D///      x137y109     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2523_1 ( .OUT(na2523_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1513_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2523_2 ( .OUT(na2523_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2523_1_i) );
// C_///AND/D      x136y107     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2524_4 ( .OUT(na2524_2_i), .IN1(na1514_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2524_5 ( .OUT(na2524_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2524_2_i) );
// C_AND/D///      x115y113     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2525_1 ( .OUT(na2525_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1515_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2525_2 ( .OUT(na2525_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2525_1_i) );
// C_///AND/D      x128y101     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2526_4 ( .OUT(na2526_2_i), .IN1(1'b1), .IN2(na1516_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2526_5 ( .OUT(na2526_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2526_2_i) );
// C_AND/D///      x106y74     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2527_1 ( .OUT(na2527_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1517_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2527_2 ( .OUT(na2527_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2527_1_i) );
// C_///AND/D      x111y102     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2528_4 ( .OUT(na2528_2_i), .IN1(na1518_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2528_5 ( .OUT(na2528_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2528_2_i) );
// C_AND/D///      x89y79     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2529_1 ( .OUT(na2529_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1519_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2529_2 ( .OUT(na2529_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2529_1_i) );
// C_///AND/D      x129y105     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2530_4 ( .OUT(na2530_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1520_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2530_5 ( .OUT(na2530_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2530_2_i) );
// C_AND/D///      x137y102     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2531_1 ( .OUT(na2531_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1521_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2531_2 ( .OUT(na2531_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2531_1_i) );
// C_///AND/D      x113y112     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2532_4 ( .OUT(na2532_2_i), .IN1(1'b1), .IN2(na1522_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2532_5 ( .OUT(na2532_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2532_2_i) );
// C_AND/D///      x115y115     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2533_1 ( .OUT(na2533_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1523_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2533_2 ( .OUT(na2533_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2533_1_i) );
// C_///AND/D      x113y90     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2534_4 ( .OUT(na2534_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1524_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2534_5 ( .OUT(na2534_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2534_2_i) );
// C_///AND/D      x99y67     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2535_4 ( .OUT(na2535_2_i), .IN1(1'b1), .IN2(na1525_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2535_5 ( .OUT(na2535_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2535_2_i) );
// C_///AND/D      x115y79     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2536_4 ( .OUT(na2536_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2536_5 ( .OUT(na2536_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2536_2_i) );
// C_AND/D///      x89y88     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2537_1 ( .OUT(na2537_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1527_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2537_2 ( .OUT(na2537_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2537_1_i) );
// C_///AND/D      x95y115     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2538_4 ( .OUT(na2538_2_i), .IN1(1'b1), .IN2(na1528_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2538_5 ( .OUT(na2538_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2538_2_i) );
// C_AND/D///      x126y107     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2539_1 ( .OUT(na2539_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1529_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2539_2 ( .OUT(na2539_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2539_1_i) );
// C_///AND/D      x110y116     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2540_4 ( .OUT(na2540_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1530_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2540_5 ( .OUT(na2540_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2540_2_i) );
// C_AND/D///      x95y116     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2541_1 ( .OUT(na2541_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1531_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2541_2 ( .OUT(na2541_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2541_1_i) );
// C_///AND/D      x94y113     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2542_4 ( .OUT(na2542_2_i), .IN1(1'b1), .IN2(na1532_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2542_5 ( .OUT(na2542_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2542_2_i) );
// C_AND/D///      x85y99     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2543_1 ( .OUT(na2543_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1533_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2543_2 ( .OUT(na2543_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2543_1_i) );
// C_///AND/D      x88y99     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2544_4 ( .OUT(na2544_2_i), .IN1(1'b1), .IN2(na1534_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2544_5 ( .OUT(na2544_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2544_2_i) );
// C_AND/D///      x85y98     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2545_1 ( .OUT(na2545_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1535_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2545_2 ( .OUT(na2545_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2545_1_i) );
// C_///AND/D      x89y105     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2546_4 ( .OUT(na2546_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1536_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2546_5 ( .OUT(na2546_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2546_2_i) );
// C_AND/D///      x99y108     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2547_1 ( .OUT(na2547_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1537_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2547_2 ( .OUT(na2547_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2547_1_i) );
// C_///AND/D      x86y80     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2548_4 ( .OUT(na2548_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1538_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2548_5 ( .OUT(na2548_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2548_2_i) );
// C_AND/D///      x91y115     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2549_1 ( .OUT(na2549_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1539_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2549_2 ( .OUT(na2549_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2549_1_i) );
// C_///AND/D      x85y76     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2550_4 ( .OUT(na2550_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1540_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2550_5 ( .OUT(na2550_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2550_2_i) );
// C_AND/D///      x88y85     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2551_1 ( .OUT(na2551_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1541_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2551_2 ( .OUT(na2551_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2551_1_i) );
// C_///AND/D      x91y79     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2552_4 ( .OUT(na2552_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1542_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2552_5 ( .OUT(na2552_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2552_2_i) );
// C_AND/D///      x89y69     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2553_1 ( .OUT(na2553_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1543_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2553_2 ( .OUT(na2553_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2553_1_i) );
// C_///AND/D      x113y116     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2554_4 ( .OUT(na2554_2_i), .IN1(1'b1), .IN2(na1544_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2554_5 ( .OUT(na2554_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2554_2_i) );
// C_AND/D///      x137y106     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2555_1 ( .OUT(na2555_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1545_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2555_2 ( .OUT(na2555_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2555_1_i) );
// C_///AND/D      x133y106     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2556_4 ( .OUT(na2556_2_i), .IN1(1'b1), .IN2(na1546_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2556_5 ( .OUT(na2556_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2556_2_i) );
// C_AND/D///      x107y115     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2557_1 ( .OUT(na2557_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1547_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2557_2 ( .OUT(na2557_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2557_1_i) );
// C_///AND/D      x124y95     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2558_4 ( .OUT(na2558_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1548_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2558_5 ( .OUT(na2558_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2558_2_i) );
// C_AND/D///      x105y73     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2559_1 ( .OUT(na2559_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1549_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2559_2 ( .OUT(na2559_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2559_1_i) );
// C_///AND/D      x115y99     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2560_4 ( .OUT(na2560_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1550_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2560_5 ( .OUT(na2560_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2560_2_i) );
// C_AND/D///      x90y79     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2561_1 ( .OUT(na2561_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1551_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2561_2 ( .OUT(na2561_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2561_1_i) );
// C_///AND/D      x132y105     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2562_4 ( .OUT(na2562_2_i), .IN1(1'b1), .IN2(na1552_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2562_5 ( .OUT(na2562_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2562_2_i) );
// C_AND/D///      x137y101     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2563_1 ( .OUT(na2563_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1553_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2563_2 ( .OUT(na2563_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2563_1_i) );
// C_AND/D///      x115y111     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2564_1 ( .OUT(na2564_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1554_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2564_2 ( .OUT(na2564_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2564_1_i) );
// C_AND/D///      x116y116     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2565_1 ( .OUT(na2565_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1555_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2565_2 ( .OUT(na2565_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2565_1_i) );
// C_///AND/D      x109y85     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2566_4 ( .OUT(na2566_2_i), .IN1(na1556_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2566_5 ( .OUT(na2566_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2566_2_i) );
// C_AND/D///      x101y67     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2567_1 ( .OUT(na2567_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1557_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2567_2 ( .OUT(na2567_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2567_1_i) );
// C_///AND/D      x119y77     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2568_4 ( .OUT(na2568_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1558_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2568_5 ( .OUT(na2568_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2568_2_i) );
// C_AND/D///      x87y87     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2569_1 ( .OUT(na2569_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1559_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2569_2 ( .OUT(na2569_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2569_1_i) );
// C_///AND/D      x95y117     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2570_4 ( .OUT(na2570_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1560_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2570_5 ( .OUT(na2570_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2570_2_i) );
// C_AND/D///      x129y108     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2571_1 ( .OUT(na2571_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1561_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2571_2 ( .OUT(na2571_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2571_1_i) );
// C_///AND/D      x107y115     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2572_4 ( .OUT(na2572_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1562_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2572_5 ( .OUT(na2572_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2572_2_i) );
// C_AND/D///      x99y117     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2573_1 ( .OUT(na2573_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1563_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2573_2 ( .OUT(na2573_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2573_1_i) );
// C_///AND/D      x87y108     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2574_4 ( .OUT(na2574_2_i), .IN1(na1564_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2574_5 ( .OUT(na2574_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2574_2_i) );
// C_AND/D///      x87y95     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2575_1 ( .OUT(na2575_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1565_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2575_2 ( .OUT(na2575_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2575_1_i) );
// C_///AND/D      x88y100     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2576_4 ( .OUT(na2576_2_i), .IN1(1'b1), .IN2(na1566_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2576_5 ( .OUT(na2576_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2576_2_i) );
// C_AND/D///      x87y96     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2577_1 ( .OUT(na2577_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1567_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2577_2 ( .OUT(na2577_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2577_1_i) );
// C_///AND/D      x85y103     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2578_4 ( .OUT(na2578_2_i), .IN1(1'b1), .IN2(na1568_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2578_5 ( .OUT(na2578_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2578_2_i) );
// C_AND/D///      x99y110     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2579_1 ( .OUT(na2579_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1569_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2579_2 ( .OUT(na2579_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2579_1_i) );
// C_///AND/D      x99y69     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2580_4 ( .OUT(na2580_2_i), .IN1(na1570_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2580_5 ( .OUT(na2580_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2580_2_i) );
// C_AND/D///      x93y113     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2581_1 ( .OUT(na2581_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1571_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2581_2 ( .OUT(na2581_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2581_1_i) );
// C_///AND/D      x93y72     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2582_4 ( .OUT(na2582_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1572_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2582_5 ( .OUT(na2582_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2582_2_i) );
// C_AND/D///      x91y85     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2583_1 ( .OUT(na2583_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1573_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2583_2 ( .OUT(na2583_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2583_1_i) );
// C_///AND/D      x89y83     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2584_4 ( .OUT(na2584_2_i), .IN1(1'b1), .IN2(na1574_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2584_5 ( .OUT(na2584_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2584_2_i) );
// C_AND/D///      x93y69     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2585_1 ( .OUT(na2585_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1575_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2585_2 ( .OUT(na2585_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2585_1_i) );
// C_///AND/D      x111y115     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2586_4 ( .OUT(na2586_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1576_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2586_5 ( .OUT(na2586_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2586_2_i) );
// C_AND/D///      x133y106     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2587_1 ( .OUT(na2587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1577_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2587_2 ( .OUT(na2587_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2587_1_i) );
// C_///AND/D      x128y99     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2588_4 ( .OUT(na2588_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1578_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2588_5 ( .OUT(na2588_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2588_2_i) );
// C_AND/D///      x103y113     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2589_1 ( .OUT(na2589_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1579_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2589_2 ( .OUT(na2589_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2589_1_i) );
// C_///AND/D      x113y93     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2590_4 ( .OUT(na2590_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1580_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2590_5 ( .OUT(na2590_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2590_2_i) );
// C_AND/D///      x101y76     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2591_1 ( .OUT(na2591_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1581_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2591_2 ( .OUT(na2591_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2591_1_i) );
// C_///AND/D      x117y103     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2592_4 ( .OUT(na2592_2_i), .IN1(na1582_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2592_5 ( .OUT(na2592_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2592_2_i) );
// C_AND/D///      x91y73     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2593_1 ( .OUT(na2593_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1583_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2593_2 ( .OUT(na2593_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2593_1_i) );
// C_AND/D///      x127y105     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2594_1 ( .OUT(na2594_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1584_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2594_2 ( .OUT(na2594_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2594_1_i) );
// C_AND/D///      x136y101     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2595_1 ( .OUT(na2595_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1585_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2595_2 ( .OUT(na2595_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2595_1_i) );
// C_///AND/D      x115y111     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2596_4 ( .OUT(na2596_2_i), .IN1(1'b1), .IN2(na1586_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2596_5 ( .OUT(na2596_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2596_2_i) );
// C_AND/D///      x119y113     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2597_1 ( .OUT(na2597_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1587_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2597_2 ( .OUT(na2597_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2597_1_i) );
// C_///AND/D      x106y89     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2598_4 ( .OUT(na2598_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1588_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2598_5 ( .OUT(na2598_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2598_2_i) );
// C_AND/D///      x105y68     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2599_1 ( .OUT(na2599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1589_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2599_2 ( .OUT(na2599_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2599_1_i) );
// C_///AND/D      x114y80     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2600_4 ( .OUT(na2600_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1590_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2600_5 ( .OUT(na2600_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2600_2_i) );
// C_AND/D///      x89y83     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2601_1 ( .OUT(na2601_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1591_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2601_2 ( .OUT(na2601_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2601_1_i) );
// C_///AND/D      x98y114     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2602_4 ( .OUT(na2602_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1592_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2602_5 ( .OUT(na2602_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2602_2_i) );
// C_AND/D///      x127y107     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2603_1 ( .OUT(na2603_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1593_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2603_2 ( .OUT(na2603_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2603_1_i) );
// C_///AND/D      x111y113     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2604_4 ( .OUT(na2604_2_i), .IN1(na1594_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2604_5 ( .OUT(na2604_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2604_2_i) );
// C_AND/D///      x98y115     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2605_1 ( .OUT(na2605_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1595_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2605_2 ( .OUT(na2605_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2605_1_i) );
// C_///AND/D      x94y109     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2606_4 ( .OUT(na2606_2_i), .IN1(na1596_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2606_5 ( .OUT(na2606_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2606_2_i) );
// C_AND/D///      x94y95     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2607_1 ( .OUT(na2607_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1597_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2607_2 ( .OUT(na2607_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2607_1_i) );
// C_///AND/D      x89y93     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2608_4 ( .OUT(na2608_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1598_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2608_5 ( .OUT(na2608_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2608_2_i) );
// C_AND/D///      x90y95     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2609_1 ( .OUT(na2609_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1599_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2609_2 ( .OUT(na2609_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2609_1_i) );
// C_///AND/D      x87y101     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2610_4 ( .OUT(na2610_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1600_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2610_5 ( .OUT(na2610_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2610_2_i) );
// C_AND/D///      x113y112     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2611_1 ( .OUT(na2611_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1601_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2611_2 ( .OUT(na2611_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2611_1_i) );
// C_///AND/D      x100y75     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2612_4 ( .OUT(na2612_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1602_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2612_5 ( .OUT(na2612_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2612_2_i) );
// C_AND/D///      x93y116     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2613_1 ( .OUT(na2613_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1603_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2613_2 ( .OUT(na2613_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2613_1_i) );
// C_///AND/D      x87y87     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2614_4 ( .OUT(na2614_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1604_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2614_5 ( .OUT(na2614_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2614_2_i) );
// C_AND/D///      x103y85     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2615_1 ( .OUT(na2615_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1605_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2615_2 ( .OUT(na2615_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2615_1_i) );
// C_///AND/D      x93y89     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2616_4 ( .OUT(na2616_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1606_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2616_5 ( .OUT(na2616_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2616_2_i) );
// C_AND/D///      x101y69     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2617_1 ( .OUT(na2617_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1607_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2617_2 ( .OUT(na2617_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2617_1_i) );
// C_///AND/D      x116y113     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2618_4 ( .OUT(na2618_2_i), .IN1(1'b1), .IN2(na1608_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2618_5 ( .OUT(na2618_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2618_2_i) );
// C_AND/D///      x135y101     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2619_1 ( .OUT(na2619_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1609_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2619_2 ( .OUT(na2619_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2619_1_i) );
// C_///AND/D      x132y109     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2620_4 ( .OUT(na2620_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1610_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2620_5 ( .OUT(na2620_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2620_2_i) );
// C_AND/D///      x112y111     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2621_1 ( .OUT(na2621_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1611_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2621_2 ( .OUT(na2621_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2621_1_i) );
// C_///AND/D      x123y92     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2622_4 ( .OUT(na2622_2_i), .IN1(na1612_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2622_5 ( .OUT(na2622_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2622_2_i) );
// C_///AND/D      x101y67     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2623_4 ( .OUT(na2623_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1613_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2623_5 ( .OUT(na2623_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2623_2_i) );
// C_///AND/D      x113y104     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2624_4 ( .OUT(na2624_2_i), .IN1(1'b1), .IN2(na1614_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2624_5 ( .OUT(na2624_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2624_2_i) );
// C_AND/D///      x100y67     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2625_1 ( .OUT(na2625_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1615_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2625_2 ( .OUT(na2625_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2625_1_i) );
// C_///AND/D      x127y101     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2626_4 ( .OUT(na2626_2_i), .IN1(1'b1), .IN2(na1616_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2626_5 ( .OUT(na2626_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2626_2_i) );
// C_AND/D///      x141y105     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2627_1 ( .OUT(na2627_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1617_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2627_2 ( .OUT(na2627_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2627_1_i) );
// C_///AND/D      x119y111     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2628_4 ( .OUT(na2628_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1618_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2628_5 ( .OUT(na2628_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2628_2_i) );
// C_AND/D///      x122y110     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2629_1 ( .OUT(na2629_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1619_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2629_2 ( .OUT(na2629_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2629_1_i) );
// C_///AND/D      x105y73     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2630_4 ( .OUT(na2630_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1620_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2630_5 ( .OUT(na2630_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2630_2_i) );
// C_AND/D///      x105y67     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2631_1 ( .OUT(na2631_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1621_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2631_2 ( .OUT(na2631_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2631_1_i) );
// C_///AND/D      x119y84     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2632_4 ( .OUT(na2632_2_i), .IN1(1'b1), .IN2(na1622_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2632_5 ( .OUT(na2632_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2632_2_i) );
// C_AND/D///      x98y84     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2633_1 ( .OUT(na2633_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1623_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2633_2 ( .OUT(na2633_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2633_1_i) );
// C_///AND/D      x95y118     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2634_4 ( .OUT(na2634_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1624_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2634_5 ( .OUT(na2634_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2634_2_i) );
// C_AND/D///      x132y107     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2635_1 ( .OUT(na2635_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1625_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2635_2 ( .OUT(na2635_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2635_1_i) );
// C_///AND/D      x109y116     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2636_4 ( .OUT(na2636_2_i), .IN1(1'b1), .IN2(na1626_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2636_5 ( .OUT(na2636_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2636_2_i) );
// C_AND/D///      x111y115     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2637_1 ( .OUT(na2637_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1627_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2637_2 ( .OUT(na2637_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2637_1_i) );
// C_///AND/D      x99y108     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2638_4 ( .OUT(na2638_2_i), .IN1(na1628_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2638_5 ( .OUT(na2638_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2638_2_i) );
// C_AND/D///      x104y83     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2639_1 ( .OUT(na2639_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1629_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2639_2 ( .OUT(na2639_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2639_1_i) );
// C_///AND/D      x97y97     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2640_4 ( .OUT(na2640_2_i), .IN1(1'b1), .IN2(na1630_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2640_5 ( .OUT(na2640_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2640_2_i) );
// C_AND/D///      x93y93     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2641_1 ( .OUT(na2641_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1631_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2641_2 ( .OUT(na2641_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2641_1_i) );
// C_///AND/D      x87y109     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2642_4 ( .OUT(na2642_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1632_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2642_5 ( .OUT(na2642_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2642_2_i) );
// C_AND/D///      x107y109     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2643_1 ( .OUT(na2643_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1633_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2643_2 ( .OUT(na2643_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2643_1_i) );
// C_///AND/D      x89y79     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2644_4 ( .OUT(na2644_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1634_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2644_5 ( .OUT(na2644_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2644_2_i) );
// C_AND/D///      x90y115     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2645_1 ( .OUT(na2645_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1635_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2645_2 ( .OUT(na2645_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2645_1_i) );
// C_///AND/D      x87y88     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2646_4 ( .OUT(na2646_2_i), .IN1(na1636_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2646_5 ( .OUT(na2646_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2646_2_i) );
// C_AND/D///      x93y79     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2647_1 ( .OUT(na2647_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1637_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2647_2 ( .OUT(na2647_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2647_1_i) );
// C_///AND/D      x89y88     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2648_4 ( .OUT(na2648_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1638_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2648_5 ( .OUT(na2648_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2648_2_i) );
// C_AND/D///      x97y70     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2649_1 ( .OUT(na2649_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1639_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2649_2 ( .OUT(na2649_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2649_1_i) );
// C_///AND/D      x109y118     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2650_4 ( .OUT(na2650_2_i), .IN1(na1640_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2650_5 ( .OUT(na2650_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2650_2_i) );
// C_AND/D///      x138y106     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2651_1 ( .OUT(na2651_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1641_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2651_2 ( .OUT(na2651_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2651_1_i) );
// C_///AND/D      x124y108     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2652_4 ( .OUT(na2652_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1642_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2652_5 ( .OUT(na2652_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2652_2_i) );
// C_///AND/D      x117y113     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2653_4 ( .OUT(na2653_2_i), .IN1(na1643_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2653_5 ( .OUT(na2653_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2653_2_i) );
// C_///AND/D      x127y105     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2654_4 ( .OUT(na2654_2_i), .IN1(1'b1), .IN2(na1644_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2654_5 ( .OUT(na2654_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2654_2_i) );
// C_AND/D///      x107y67     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2655_1 ( .OUT(na2655_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1645_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2655_2 ( .OUT(na2655_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2655_1_i) );
// C_///AND/D      x100y107     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2656_4 ( .OUT(na2656_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1646_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2656_5 ( .OUT(na2656_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2656_2_i) );
// C_AND/D///      x93y67     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2657_1 ( .OUT(na2657_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1647_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2657_2 ( .OUT(na2657_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2657_1_i) );
// C_///AND/D      x126y107     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2658_4 ( .OUT(na2658_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1648_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2658_5 ( .OUT(na2658_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2658_2_i) );
// C_AND/D///      x133y102     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2659_1 ( .OUT(na2659_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1649_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2659_2 ( .OUT(na2659_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2659_1_i) );
// C_///AND/D      x115y113     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2660_4 ( .OUT(na2660_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1650_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2660_5 ( .OUT(na2660_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2660_2_i) );
// C_AND/D///      x117y113     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2661_1 ( .OUT(na2661_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1651_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2661_2 ( .OUT(na2661_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2661_1_i) );
// C_///AND/D      x113y91     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2662_4 ( .OUT(na2662_2_i), .IN1(1'b1), .IN2(na1652_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2662_5 ( .OUT(na2662_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2662_2_i) );
// C_AND/D///      x103y68     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2663_1 ( .OUT(na2663_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1653_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2663_2 ( .OUT(na2663_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2663_1_i) );
// C_///AND/D      x116y87     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2664_4 ( .OUT(na2664_2_i), .IN1(na1654_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2664_5 ( .OUT(na2664_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2664_2_i) );
// C_AND/D///      x87y81     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2665_1 ( .OUT(na2665_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1655_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2665_2 ( .OUT(na2665_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2665_1_i) );
// C_///AND/D      x93y116     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2666_4 ( .OUT(na2666_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1656_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2666_5 ( .OUT(na2666_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2666_2_i) );
// C_AND/D///      x132y105     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2667_1 ( .OUT(na2667_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1657_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2667_2 ( .OUT(na2667_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2667_1_i) );
// C_///AND/D      x104y117     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2668_4 ( .OUT(na2668_2_i), .IN1(na1658_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2668_5 ( .OUT(na2668_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2668_2_i) );
// C_AND/D///      x101y116     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2669_1 ( .OUT(na2669_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1659_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2669_2 ( .OUT(na2669_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2669_1_i) );
// C_///AND/D      x91y107     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2670_4 ( .OUT(na2670_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1660_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2670_5 ( .OUT(na2670_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2670_2_i) );
// C_AND/D///      x95y91     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2671_1 ( .OUT(na2671_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1661_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2671_2 ( .OUT(na2671_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2671_1_i) );
// C_///AND/D      x94y105     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2672_4 ( .OUT(na2672_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1662_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2672_5 ( .OUT(na2672_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2672_2_i) );
// C_AND/D///      x87y93     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2673_1 ( .OUT(na2673_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1663_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2673_2 ( .OUT(na2673_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2673_1_i) );
// C_///AND/D      x85y108     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2674_4 ( .OUT(na2674_2_i), .IN1(na1664_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2674_5 ( .OUT(na2674_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2674_2_i) );
// C_AND/D///      x104y110     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2675_1 ( .OUT(na2675_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1665_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2675_2 ( .OUT(na2675_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2675_1_i) );
// C_///AND/D      x92y77     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2676_4 ( .OUT(na2676_2_i), .IN1(na1666_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2676_5 ( .OUT(na2676_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2676_2_i) );
// C_AND/D///      x92y115     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2677_1 ( .OUT(na2677_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1667_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2677_2 ( .OUT(na2677_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2677_1_i) );
// C_///AND/D      x87y84     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2678_4 ( .OUT(na2678_2_i), .IN1(na1668_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2678_5 ( .OUT(na2678_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2678_2_i) );
// C_AND/D///      x91y79     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2679_1 ( .OUT(na2679_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1669_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2679_2 ( .OUT(na2679_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2679_1_i) );
// C_///AND/D      x93y92     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2680_4 ( .OUT(na2680_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1670_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2680_5 ( .OUT(na2680_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2680_2_i) );
// C_AND/D///      x94y68     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2681_1 ( .OUT(na2681_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1671_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2681_2 ( .OUT(na2681_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2681_1_i) );
// C_AND/D///      x109y115     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2682_1 ( .OUT(na2682_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1672_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2682_2 ( .OUT(na2682_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2682_1_i) );
// C_AND/D///      x139y106     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2683_1 ( .OUT(na2683_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1673_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2683_2 ( .OUT(na2683_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2683_1_i) );
// C_///AND/D      x127y111     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2684_4 ( .OUT(na2684_2_i), .IN1(1'b1), .IN2(na1674_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2684_5 ( .OUT(na2684_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2684_2_i) );
// C_AND/D///      x111y113     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2685_1 ( .OUT(na2685_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1675_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2685_2 ( .OUT(na2685_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2685_1_i) );
// C_///AND/D      x121y102     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2686_4 ( .OUT(na2686_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1676_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2686_5 ( .OUT(na2686_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2686_2_i) );
// C_AND/D///      x104y70     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2687_1 ( .OUT(na2687_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1677_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2687_2 ( .OUT(na2687_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2687_1_i) );
// C_///AND/D      x109y105     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2688_4 ( .OUT(na2688_2_i), .IN1(na1678_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2688_5 ( .OUT(na2688_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2688_2_i) );
// C_AND/D///      x93y65     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2689_1 ( .OUT(na2689_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1679_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2689_2 ( .OUT(na2689_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2689_1_i) );
// C_///AND/D      x131y107     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2690_4 ( .OUT(na2690_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1680_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2690_5 ( .OUT(na2690_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2690_2_i) );
// C_AND/D///      x139y101     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2691_1 ( .OUT(na2691_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1681_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2691_2 ( .OUT(na2691_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2691_1_i) );
// C_///AND/D      x115y112     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2692_4 ( .OUT(na2692_2_i), .IN1(na1682_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2692_5 ( .OUT(na2692_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2692_2_i) );
// C_AND/D///      x116y114     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2693_1 ( .OUT(na2693_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1683_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2693_2 ( .OUT(na2693_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2693_1_i) );
// C_///AND/D      x109y88     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2694_4 ( .OUT(na2694_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1684_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2694_5 ( .OUT(na2694_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2694_2_i) );
// C_AND/D///      x100y66     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2695_1 ( .OUT(na2695_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1685_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2695_2 ( .OUT(na2695_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2695_1_i) );
// C_///AND/D      x116y81     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2696_4 ( .OUT(na2696_2_i), .IN1(na1686_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2696_5 ( .OUT(na2696_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2696_2_i) );
// C_AND/D///      x87y84     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2697_1 ( .OUT(na2697_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1687_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2697_2 ( .OUT(na2697_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2697_1_i) );
// C_///AND/D      x93y113     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2698_4 ( .OUT(na2698_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1688_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2698_5 ( .OUT(na2698_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2698_2_i) );
// C_AND/D///      x132y108     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2699_1 ( .OUT(na2699_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1689_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2699_2 ( .OUT(na2699_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2699_1_i) );
// C_///AND/D      x107y118     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2700_4 ( .OUT(na2700_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1690_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2700_5 ( .OUT(na2700_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2700_2_i) );
// C_AND/D///      x102y116     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2701_1 ( .OUT(na2701_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1691_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2701_2 ( .OUT(na2701_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2701_1_i) );
// C_///AND/D      x93y106     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2702_4 ( .OUT(na2702_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1692_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2702_5 ( .OUT(na2702_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2702_2_i) );
// C_AND/D///      x93y89     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2703_1 ( .OUT(na2703_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1693_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2703_2 ( .OUT(na2703_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2703_1_i) );
// C_///AND/D      x93y104     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2704_4 ( .OUT(na2704_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1694_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2704_5 ( .OUT(na2704_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2704_2_i) );
// C_AND/D///      x89y93     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2705_1 ( .OUT(na2705_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1695_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2705_2 ( .OUT(na2705_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2705_1_i) );
// C_///AND/D      x87y106     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2706_4 ( .OUT(na2706_2_i), .IN1(1'b1), .IN2(na1696_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2706_5 ( .OUT(na2706_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2706_2_i) );
// C_AND/D///      x105y108     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2707_1 ( .OUT(na2707_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1697_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2707_2 ( .OUT(na2707_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2707_1_i) );
// C_///AND/D      x101y76     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2708_4 ( .OUT(na2708_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1698_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2708_5 ( .OUT(na2708_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2708_2_i) );
// C_AND/D///      x94y115     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2709_1 ( .OUT(na2709_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1699_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2709_2 ( .OUT(na2709_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2709_1_i) );
// C_///AND/D      x89y85     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2710_4 ( .OUT(na2710_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1700_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2710_5 ( .OUT(na2710_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2710_2_i) );
// C_///AND/D      x94y71     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2711_4 ( .OUT(na2711_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1701_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2711_5 ( .OUT(na2711_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2711_2_i) );
// C_///AND/D      x93y93     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2712_4 ( .OUT(na2712_2_i), .IN1(na1702_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2712_5 ( .OUT(na2712_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2712_2_i) );
// C_AND/D///      x99y65     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2713_1 ( .OUT(na2713_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1703_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2713_2 ( .OUT(na2713_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2713_1_i) );
// C_///AND/D      x109y115     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2714_4 ( .OUT(na2714_2_i), .IN1(1'b1), .IN2(na1704_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2714_5 ( .OUT(na2714_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2714_2_i) );
// C_AND/D///      x135y105     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2715_1 ( .OUT(na2715_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1705_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2715_2 ( .OUT(na2715_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2715_1_i) );
// C_///AND/D      x123y108     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2716_4 ( .OUT(na2716_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1706_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2716_5 ( .OUT(na2716_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2716_2_i) );
// C_AND/D///      x113y113     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2717_1 ( .OUT(na2717_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1707_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2717_2 ( .OUT(na2717_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2717_1_i) );
// C_///AND/D      x121y96     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2718_4 ( .OUT(na2718_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1708_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2718_5 ( .OUT(na2718_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2718_2_i) );
// C_AND/D///      x105y72     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2719_1 ( .OUT(na2719_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1709_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2719_2 ( .OUT(na2719_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2719_1_i) );
// C_///AND/D      x109y103     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2720_4 ( .OUT(na2720_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1710_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2720_5 ( .OUT(na2720_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2720_2_i) );
// C_AND/D///      x97y65     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2721_1 ( .OUT(na2721_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1711_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2721_2 ( .OUT(na2721_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2721_1_i) );
// C_///AND/D      x127y107     80'hC0_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2722_4 ( .OUT(na2722_2_i), .IN1(1'b1), .IN2(na1712_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2722_5 ( .OUT(na2722_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2722_2_i) );
// C_AND/D///      x134y101     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2723_1 ( .OUT(na2723_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1713_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2723_2 ( .OUT(na2723_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2723_1_i) );
// C_///AND/D      x114y111     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2724_4 ( .OUT(na2724_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1714_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2724_5 ( .OUT(na2724_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2724_2_i) );
// C_AND/D///      x115y112     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2725_1 ( .OUT(na2725_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1715_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2725_2 ( .OUT(na2725_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2725_1_i) );
// C_///AND/D      x104y89     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2726_4 ( .OUT(na2726_2_i), .IN1(na1716_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2726_5 ( .OUT(na2726_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2726_2_i) );
// C_AND/D///      x99y67     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2727_1 ( .OUT(na2727_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1717_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2727_2 ( .OUT(na2727_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2727_1_i) );
// C_///AND/D      x113y83     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2728_4 ( .OUT(na2728_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1718_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2728_5 ( .OUT(na2728_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2728_2_i) );
// C_AND/D///      x91y84     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2729_1 ( .OUT(na2729_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1719_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2729_2 ( .OUT(na2729_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2729_1_i) );
// C_///AND/D      x91y116     80'hC0_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2730_4 ( .OUT(na2730_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1720_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2730_5 ( .OUT(na2730_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2730_2_i) );
// C_AND/D///      x129y105     80'hC0_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2731_1 ( .OUT(na2731_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1721_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2731_2 ( .OUT(na2731_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2731_1_i) );
// C_///AND/D      x115y116     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2732_4 ( .OUT(na2732_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1722_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2732_5 ( .OUT(na2732_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2732_2_i) );
// C_AND/D///      x106y113     80'hC0_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2733_1 ( .OUT(na2733_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1723_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2733_2 ( .OUT(na2733_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2733_1_i) );
// C_///AND/D      x91y104     80'hC0_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2734_4 ( .OUT(na2734_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1724_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2734_5 ( .OUT(na2734_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2734_2_i) );
// C_AND/D///      x95y89     80'hC0_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2735_1 ( .OUT(na2735_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1725_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2735_2 ( .OUT(na2735_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2735_1_i) );
// C_///AND/D      x93y98     80'hC0_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2736_4 ( .OUT(na2736_2_i), .IN1(na1726_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a2736_5 ( .OUT(na2736_2), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2736_2_i) );
// C_AND/D///      x92y93     80'hC0_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2737_1 ( .OUT(na2737_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1727_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a2737_2 ( .OUT(na2737_1), .CLK(1'b0), .EN(1'b0), .SR(na3277_1), .CINY2(na4481_3), .PINY2(~na4481_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2737_1_i) );
// C_///AND/D      x87y102     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2738_4 ( .OUT(na2738_2_i), .IN1(na607_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2738_5 ( .OUT(na2738_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2738_2_i) );
// C_AND/D///      x101y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2739_1 ( .OUT(na2739_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na608_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2739_2 ( .OUT(na2739_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2739_1_i) );
// C_AND/D///      x99y84     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2740_1 ( .OUT(na2740_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na609_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2740_2 ( .OUT(na2740_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2740_1_i) );
// C_AND/D///      x91y109     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2741_1 ( .OUT(na2741_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na610_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2741_2 ( .OUT(na2741_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2741_1_i) );
// C_///AND/D      x91y75     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2742_4 ( .OUT(na2742_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na611_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2742_5 ( .OUT(na2742_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2742_2_i) );
// C_AND/D///      x96y86     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2743_1 ( .OUT(na2743_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na612_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2743_2 ( .OUT(na2743_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2743_1_i) );
// C_///AND/D      x94y67     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2745_4 ( .OUT(na2745_2_i), .IN1(na614_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2745_5 ( .OUT(na2745_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2745_2_i) );
// C_AND/D///      x114y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2746_1 ( .OUT(na2746_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na615_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2746_2 ( .OUT(na2746_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2746_1_i) );
// C_///AND/D      x131y108     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2748_4 ( .OUT(na2748_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na617_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2748_5 ( .OUT(na2748_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2748_2_i) );
// C_AND/D///      x116y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2749_1 ( .OUT(na2749_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na618_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2749_2 ( .OUT(na2749_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2749_1_i) );
// C_///AND/D      x127y89     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2750_4 ( .OUT(na2750_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na619_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2750_5 ( .OUT(na2750_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2750_2_i) );
// C_AND/D///      x111y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2752_1 ( .OUT(na2752_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na621_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2752_2 ( .OUT(na2752_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2752_1_i) );
// C_///AND/D      x98y72     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2753_4 ( .OUT(na2753_2_i), .IN1(na622_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2753_5 ( .OUT(na2753_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2753_2_i) );
// C_AND/D///      x115y101     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2756_1 ( .OUT(na2756_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na625_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2756_2 ( .OUT(na2756_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2756_1_i) );
// C_///AND/D      x121y105     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2757_4 ( .OUT(na2757_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na626_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2757_5 ( .OUT(na2757_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2757_2_i) );
// C_AND/D///      x115y85     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2758_1 ( .OUT(na2758_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na627_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2758_2 ( .OUT(na2758_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2758_1_i) );
// C_///AND/D      x103y65     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2759_4 ( .OUT(na2759_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na628_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2759_5 ( .OUT(na2759_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2759_2_i) );
// C_AND/D///      x100y85     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2761_1 ( .OUT(na2761_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na630_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2761_2 ( .OUT(na2761_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2761_1_i) );
// C_///AND/D      x96y111     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2762_4 ( .OUT(na2762_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na631_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2762_5 ( .OUT(na2762_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2762_2_i) );
// C_AND/D///      x125y108     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2763_1 ( .OUT(na2763_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na632_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2763_2 ( .OUT(na2763_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2763_1_i) );
// C_///AND/D      x112y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2764_4 ( .OUT(na2764_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na633_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2764_5 ( .OUT(na2764_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2764_2_i) );
// C_AND/D///      x104y111     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2765_1 ( .OUT(na2765_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na634_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2765_2 ( .OUT(na2765_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2765_1_i) );
// C_///AND/D      x93y108     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2766_4 ( .OUT(na2766_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na635_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2766_5 ( .OUT(na2766_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2766_2_i) );
// C_AND/D///      x91y98     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2767_1 ( .OUT(na2767_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na636_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2767_2 ( .OUT(na2767_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2767_1_i) );
// C_///AND/D      x89y104     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2768_4 ( .OUT(na2768_2_i), .IN1(1'b1), .IN2(na637_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2768_5 ( .OUT(na2768_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2768_2_i) );
// C_AND/D///      x95y101     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2769_1 ( .OUT(na2769_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na638_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2769_2 ( .OUT(na2769_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2769_1_i) );
// C_///AND/D      x87y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2770_4 ( .OUT(na2770_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na639_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2770_5 ( .OUT(na2770_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2770_2_i) );
// C_AND/D///      x105y105     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2771_1 ( .OUT(na2771_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na640_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2771_2 ( .OUT(na2771_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2771_1_i) );
// C_///AND/D      x100y71     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2772_4 ( .OUT(na2772_2_i), .IN1(na641_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2772_5 ( .OUT(na2772_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2772_2_i) );
// C_AND/D///      x87y114     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2773_1 ( .OUT(na2773_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na642_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2773_2 ( .OUT(na2773_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2773_1_i) );
// C_///AND/D      x88y78     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2774_4 ( .OUT(na2774_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na643_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2774_5 ( .OUT(na2774_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2774_2_i) );
// C_AND/D///      x91y87     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2775_1 ( .OUT(na2775_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na644_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2775_2 ( .OUT(na2775_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2775_1_i) );
// C_AND/D///      x94y87     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2776_1 ( .OUT(na2776_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na645_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2776_2 ( .OUT(na2776_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2776_1_i) );
// C_AND/D///      x98y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2777_1 ( .OUT(na2777_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na646_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2777_2 ( .OUT(na2777_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2777_1_i) );
// C_///AND/D      x117y115     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2778_4 ( .OUT(na2778_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na647_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2778_5 ( .OUT(na2778_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2778_2_i) );
// C_AND/D///      x137y104     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2779_1 ( .OUT(na2779_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na648_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2779_2 ( .OUT(na2779_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2779_1_i) );
// C_///AND/D      x139y105     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2780_4 ( .OUT(na2780_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na649_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2780_5 ( .OUT(na2780_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2780_2_i) );
// C_AND/D///      x111y111     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2781_1 ( .OUT(na2781_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na650_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2781_2 ( .OUT(na2781_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2781_1_i) );
// C_///AND/D      x123y100     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2782_4 ( .OUT(na2782_2_i), .IN1(1'b1), .IN2(na651_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2782_5 ( .OUT(na2782_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2782_2_i) );
// C_AND/D///      x106y73     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2783_1 ( .OUT(na2783_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na652_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2783_2 ( .OUT(na2783_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2783_1_i) );
// C_///AND/D      x113y102     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2784_4 ( .OUT(na2784_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na653_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2784_5 ( .OUT(na2784_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2784_2_i) );
// C_AND/D///      x91y75     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2785_1 ( .OUT(na2785_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na654_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2785_2 ( .OUT(na2785_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2785_1_i) );
// C_///AND/D      x133y107     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2786_4 ( .OUT(na2786_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na655_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2786_5 ( .OUT(na2786_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2786_2_i) );
// C_AND/D///      x139y100     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2787_1 ( .OUT(na2787_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na656_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2787_2 ( .OUT(na2787_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2787_1_i) );
// C_///AND/D      x121y111     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2788_4 ( .OUT(na2788_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na657_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2788_5 ( .OUT(na2788_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2788_2_i) );
// C_AND/D///      x120y115     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2789_1 ( .OUT(na2789_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na658_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2789_2 ( .OUT(na2789_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2789_1_i) );
// C_///AND/D      x117y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2790_4 ( .OUT(na2790_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na659_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2790_5 ( .OUT(na2790_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2790_2_i) );
// C_AND/D///      x105y70     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2791_1 ( .OUT(na2791_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na660_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2791_2 ( .OUT(na2791_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2791_1_i) );
// C_///AND/D      x123y77     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2792_4 ( .OUT(na2792_2_i), .IN1(1'b1), .IN2(na661_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2792_5 ( .OUT(na2792_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2792_2_i) );
// C_AND/D///      x90y88     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2793_1 ( .OUT(na2793_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na662_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2793_2 ( .OUT(na2793_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2793_1_i) );
// C_///AND/D      x94y114     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2794_4 ( .OUT(na2794_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na663_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2794_5 ( .OUT(na2794_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2794_2_i) );
// C_AND/D///      x128y108     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2795_1 ( .OUT(na2795_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na664_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2795_2 ( .OUT(na2795_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2795_1_i) );
// C_///AND/D      x111y114     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2796_4 ( .OUT(na2796_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na665_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2796_5 ( .OUT(na2796_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2796_2_i) );
// C_AND/D///      x100y116     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2797_1 ( .OUT(na2797_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na666_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2797_2 ( .OUT(na2797_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2797_1_i) );
// C_///AND/D      x95y109     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2798_4 ( .OUT(na2798_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na667_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2798_5 ( .OUT(na2798_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2798_2_i) );
// C_AND/D///      x87y97     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2799_1 ( .OUT(na2799_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na668_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2799_2 ( .OUT(na2799_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2799_1_i) );
// C_///AND/D      x92y105     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2800_4 ( .OUT(na2800_2_i), .IN1(1'b1), .IN2(na669_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2800_5 ( .OUT(na2800_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2800_2_i) );
// C_AND/D///      x86y97     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2801_1 ( .OUT(na2801_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na670_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2801_2 ( .OUT(na2801_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2801_1_i) );
// C_///AND/D      x88y102     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2802_4 ( .OUT(na2802_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na671_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2802_5 ( .OUT(na2802_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2802_2_i) );
// C_AND/D///      x103y106     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2803_1 ( .OUT(na2803_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na672_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2803_2 ( .OUT(na2803_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2803_1_i) );
// C_///AND/D      x98y74     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2804_4 ( .OUT(na2804_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na673_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2804_5 ( .OUT(na2804_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2804_2_i) );
// C_///AND/D      x92y112     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2805_4 ( .OUT(na2805_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na674_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2805_5 ( .OUT(na2805_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2805_2_i) );
// C_///AND/D      x90y71     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2806_4 ( .OUT(na2806_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na675_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2806_5 ( .OUT(na2806_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2806_2_i) );
// C_AND/D///      x94y84     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2807_1 ( .OUT(na2807_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na676_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2807_2 ( .OUT(na2807_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2807_1_i) );
// C_///AND/D      x95y80     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2808_4 ( .OUT(na2808_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na677_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2808_5 ( .OUT(na2808_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2808_2_i) );
// C_AND/D///      x96y68     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2809_1 ( .OUT(na2809_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na678_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2809_2 ( .OUT(na2809_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2809_1_i) );
// C_///AND/D      x117y114     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2810_4 ( .OUT(na2810_2_i), .IN1(1'b1), .IN2(na679_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2810_5 ( .OUT(na2810_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2810_2_i) );
// C_AND/D///      x140y106     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2811_1 ( .OUT(na2811_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na680_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2811_2 ( .OUT(na2811_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2811_1_i) );
// C_///AND/D      x133y104     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2812_4 ( .OUT(na2812_2_i), .IN1(na681_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2812_5 ( .OUT(na2812_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2812_2_i) );
// C_AND/D///      x110y113     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2813_1 ( .OUT(na2813_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na682_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2813_2 ( .OUT(na2813_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2813_1_i) );
// C_///AND/D      x126y94     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2814_4 ( .OUT(na2814_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na683_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2814_5 ( .OUT(na2814_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2814_2_i) );
// C_AND/D///      x105y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2815_1 ( .OUT(na2815_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na684_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2815_2 ( .OUT(na2815_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2815_1_i) );
// C_///AND/D      x118y101     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2816_4 ( .OUT(na2816_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na685_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2816_5 ( .OUT(na2816_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2816_2_i) );
// C_AND/D///      x95y76     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2817_1 ( .OUT(na2817_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na686_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2817_2 ( .OUT(na2817_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2817_1_i) );
// C_///AND/D      x138y103     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2818_4 ( .OUT(na2818_2_i), .IN1(1'b1), .IN2(na687_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2818_5 ( .OUT(na2818_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2818_2_i) );
// C_AND/D///      x138y100     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2819_1 ( .OUT(na2819_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na688_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2819_2 ( .OUT(na2819_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2819_1_i) );
// C_///AND/D      x123y112     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2820_4 ( .OUT(na2820_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na689_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2820_5 ( .OUT(na2820_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2820_2_i) );
// C_AND/D///      x120y112     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2821_1 ( .OUT(na2821_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na690_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2821_2 ( .OUT(na2821_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2821_1_i) );
// C_///AND/D      x119y90     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2822_4 ( .OUT(na2822_2_i), .IN1(1'b1), .IN2(na691_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2822_5 ( .OUT(na2822_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2822_2_i) );
// C_AND/D///      x106y67     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2823_1 ( .OUT(na2823_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na692_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2823_2 ( .OUT(na2823_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2823_1_i) );
// C_///AND/D      x121y76     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2824_4 ( .OUT(na2824_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na693_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2824_5 ( .OUT(na2824_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2824_2_i) );
// C_AND/D///      x89y87     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2825_1 ( .OUT(na2825_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na694_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2825_2 ( .OUT(na2825_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2825_1_i) );
// C_///AND/D      x96y113     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2826_4 ( .OUT(na2826_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na695_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2826_5 ( .OUT(na2826_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2826_2_i) );
// C_AND/D///      x130y106     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2827_1 ( .OUT(na2827_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na696_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2827_2 ( .OUT(na2827_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2827_1_i) );
// C_///AND/D      x114y114     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2828_4 ( .OUT(na2828_2_i), .IN1(na697_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2828_5 ( .OUT(na2828_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2828_2_i) );
// C_AND/D///      x102y115     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2829_1 ( .OUT(na2829_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na698_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2829_2 ( .OUT(na2829_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2829_1_i) );
// C_///AND/D      x98y108     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2830_4 ( .OUT(na2830_2_i), .IN1(1'b1), .IN2(na699_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2830_5 ( .OUT(na2830_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2830_2_i) );
// C_AND/D///      x94y94     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2831_1 ( .OUT(na2831_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na700_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2831_2 ( .OUT(na2831_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2831_1_i) );
// C_///AND/D      x90y100     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2832_4 ( .OUT(na2832_2_i), .IN1(na701_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2832_5 ( .OUT(na2832_2), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2832_2_i) );
// C_AND/D///      x92y96     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2833_1 ( .OUT(na2833_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na702_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2833_2 ( .OUT(na2833_1), .CLK(1'b0), .EN(na1460_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2833_1_i) );
// C_///AND/D      x90y101     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2834_4 ( .OUT(na2834_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na703_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2834_5 ( .OUT(na2834_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2834_2_i) );
// C_///AND/D      x116y107     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2835_4 ( .OUT(na2835_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na704_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2835_5 ( .OUT(na2835_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2835_2_i) );
// C_///AND/D      x103y75     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2836_4 ( .OUT(na2836_2_i), .IN1(na705_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2836_5 ( .OUT(na2836_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2836_2_i) );
// C_AND/D///      x93y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2837_1 ( .OUT(na2837_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na706_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2837_2 ( .OUT(na2837_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2837_1_i) );
// C_///AND/D      x88y84     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2838_4 ( .OUT(na2838_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na707_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2838_5 ( .OUT(na2838_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2838_2_i) );
// C_AND/D///      x98y82     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2839_1 ( .OUT(na2839_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na708_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2839_2 ( .OUT(na2839_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2839_1_i) );
// C_///AND/D      x99y66     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2841_4 ( .OUT(na2841_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na710_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2841_5 ( .OUT(na2841_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2841_2_i) );
// C_AND/D///      x112y112     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2842_1 ( .OUT(na2842_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na711_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2842_2 ( .OUT(na2842_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2842_1_i) );
// C_///AND/D      x129y106     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2844_4 ( .OUT(na2844_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na713_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2844_5 ( .OUT(na2844_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2844_2_i) );
// C_AND/D///      x115y109     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2845_1 ( .OUT(na2845_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na714_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2845_2 ( .OUT(na2845_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2845_1_i) );
// C_///AND/D      x121y89     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2846_4 ( .OUT(na2846_2_i), .IN1(na715_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2846_5 ( .OUT(na2846_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2846_2_i) );
// C_AND/D///      x109y99     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2848_1 ( .OUT(na2848_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na717_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2848_2 ( .OUT(na2848_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2848_1_i) );
// C_///AND/D      x102y66     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2849_4 ( .OUT(na2849_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na718_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2849_5 ( .OUT(na2849_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2849_2_i) );
// C_AND/D///      x117y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2852_1 ( .OUT(na2852_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na721_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2852_2 ( .OUT(na2852_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2852_1_i) );
// C_///AND/D      x123y105     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2853_4 ( .OUT(na2853_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na722_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2853_5 ( .OUT(na2853_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2853_2_i) );
// C_AND/D///      x113y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2854_1 ( .OUT(na2854_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na723_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2854_2 ( .OUT(na2854_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2854_1_i) );
// C_///AND/D      x105y66     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2855_4 ( .OUT(na2855_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na724_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2855_5 ( .OUT(na2855_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2855_2_i) );
// C_AND/D///      x100y84     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2857_1 ( .OUT(na2857_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na726_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2857_2 ( .OUT(na2857_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2857_1_i) );
// C_///AND/D      x95y108     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2858_4 ( .OUT(na2858_2_i), .IN1(na727_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2858_5 ( .OUT(na2858_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2858_2_i) );
// C_AND/D///      x107y111     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2860_1 ( .OUT(na2860_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na729_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2860_2 ( .OUT(na2860_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2860_1_i) );
// C_///AND/D      x112y112     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2861_4 ( .OUT(na2861_2_i), .IN1(1'b1), .IN2(na730_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2861_5 ( .OUT(na2861_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2861_2_i) );
// C_AND/D///      x97y105     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2862_1 ( .OUT(na2862_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na731_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2862_2 ( .OUT(na2862_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2862_1_i) );
// C_///AND/D      x99y83     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2863_4 ( .OUT(na2863_2_i), .IN1(na732_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2863_5 ( .OUT(na2863_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2863_2_i) );
// C_AND/D///      x97y95     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2865_1 ( .OUT(na2865_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na734_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2865_2 ( .OUT(na2865_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2865_1_i) );
// C_///AND/D      x87y104     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2866_4 ( .OUT(na2866_2_i), .IN1(1'b1), .IN2(na767_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2866_5 ( .OUT(na2866_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2866_2_i) );
// C_AND/D///      x103y105     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2867_1 ( .OUT(na2867_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na768_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2867_2 ( .OUT(na2867_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2867_1_i) );
// C_///AND/D      x104y73     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2868_4 ( .OUT(na2868_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na769_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2868_5 ( .OUT(na2868_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2868_2_i) );
// C_AND/D///      x91y114     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2869_1 ( .OUT(na2869_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na770_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2869_2 ( .OUT(na2869_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2869_1_i) );
// C_///AND/D      x99y80     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2870_4 ( .OUT(na2870_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na771_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2870_5 ( .OUT(na2870_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2870_2_i) );
// C_AND/D///      x94y81     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2871_1 ( .OUT(na2871_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na772_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2871_2 ( .OUT(na2871_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2871_1_i) );
// C_AND/D///      x100y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2872_1 ( .OUT(na2872_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na773_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2872_2 ( .OUT(na2872_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2872_1_i) );
// C_AND/D///      x99y66     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2873_1 ( .OUT(na2873_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na774_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2873_2 ( .OUT(na2873_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2873_1_i) );
// C_///AND/D      x113y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2874_4 ( .OUT(na2874_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na775_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2874_5 ( .OUT(na2874_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2874_2_i) );
// C_AND/D///      x140y103     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2875_1 ( .OUT(na2875_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na776_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2875_2 ( .OUT(na2875_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2875_1_i) );
// C_///AND/D      x128y105     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2876_4 ( .OUT(na2876_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na777_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2876_5 ( .OUT(na2876_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2876_2_i) );
// C_AND/D///      x112y113     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2877_1 ( .OUT(na2877_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na778_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2877_2 ( .OUT(na2877_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2877_1_i) );
// C_///AND/D      x124y97     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2878_4 ( .OUT(na2878_2_i), .IN1(na779_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2878_5 ( .OUT(na2878_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2878_2_i) );
// C_AND/D///      x107y69     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2879_1 ( .OUT(na2879_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na780_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2879_2 ( .OUT(na2879_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2879_1_i) );
// C_///AND/D      x111y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2880_4 ( .OUT(na2880_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na781_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2880_5 ( .OUT(na2880_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2880_2_i) );
// C_AND/D///      x99y68     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2881_1 ( .OUT(na2881_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na782_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2881_2 ( .OUT(na2881_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2881_1_i) );
// C_///AND/D      x131y104     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2882_4 ( .OUT(na2882_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na783_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2882_5 ( .OUT(na2882_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2882_2_i) );
// C_AND/D///      x137y99     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2883_1 ( .OUT(na2883_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na784_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2883_2 ( .OUT(na2883_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2883_1_i) );
// C_///AND/D      x115y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2884_4 ( .OUT(na2884_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na785_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2884_5 ( .OUT(na2884_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2884_2_i) );
// C_AND/D///      x119y112     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2885_1 ( .OUT(na2885_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na786_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2885_2 ( .OUT(na2885_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2885_1_i) );
// C_///AND/D      x114y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2886_4 ( .OUT(na2886_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na787_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2886_5 ( .OUT(na2886_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2886_2_i) );
// C_AND/D///      x104y67     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2887_1 ( .OUT(na2887_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na788_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2887_2 ( .OUT(na2887_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2887_1_i) );
// C_///AND/D      x118y79     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2888_4 ( .OUT(na2888_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na789_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2888_5 ( .OUT(na2888_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2888_2_i) );
// C_AND/D///      x92y81     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2889_1 ( .OUT(na2889_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na790_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2889_2 ( .OUT(na2889_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2889_1_i) );
// C_///AND/D      x93y114     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2890_4 ( .OUT(na2890_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na791_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2890_5 ( .OUT(na2890_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2890_2_i) );
// C_AND/D///      x133y105     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2891_1 ( .OUT(na2891_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na792_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2891_2 ( .OUT(na2891_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2891_1_i) );
// C_///AND/D      x112y113     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2892_4 ( .OUT(na2892_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na793_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2892_5 ( .OUT(na2892_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2892_2_i) );
// C_AND/D///      x108y115     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2893_1 ( .OUT(na2893_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na794_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2893_2 ( .OUT(na2893_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2893_1_i) );
// C_///AND/D      x98y107     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2894_4 ( .OUT(na2894_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na795_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2894_5 ( .OUT(na2894_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2894_2_i) );
// C_AND/D///      x98y91     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2895_1 ( .OUT(na2895_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na796_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2895_2 ( .OUT(na2895_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2895_1_i) );
// C_///AND/D      x102y95     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2896_4 ( .OUT(na2896_2_i), .IN1(1'b1), .IN2(na797_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2896_5 ( .OUT(na2896_2), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2896_2_i) );
// C_AND/D///      x89y92     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2897_1 ( .OUT(na2897_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na798_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2897_2 ( .OUT(na2897_1), .CLK(1'b0), .EN(na1462_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2897_1_i) );
// C_///AND/D      x134y85     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2898_4 ( .OUT(na2898_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1125_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2898_5 ( .OUT(na2898_2), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2898_2_i) );
// C_AND/D///      x133y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2899_1 ( .OUT(na2899_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1127_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2899_2 ( .OUT(na2899_1), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2899_1_i) );
// C_///AND/D      x135y73     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2900_4 ( .OUT(na2900_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1128_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2900_5 ( .OUT(na2900_2), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2900_2_i) );
// C_AND/D///      x127y87     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2901_1 ( .OUT(na2901_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1129_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2901_2 ( .OUT(na2901_1), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2901_1_i) );
// C_AND/D///      x131y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2902_1 ( .OUT(na2902_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2902_2 ( .OUT(na2902_1), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2902_1_i) );
// C_AND/D///      x132y75     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2903_1 ( .OUT(na2903_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1131_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2903_2 ( .OUT(na2903_1), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2903_1_i) );
// C_///AND/D      x134y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2904_4 ( .OUT(na2904_2_i), .IN1(1'b1), .IN2(na1132_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2904_5 ( .OUT(na2904_2), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2904_2_i) );
// C_AND/D///      x131y73     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2905_1 ( .OUT(na2905_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1133_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2905_2 ( .OUT(na2905_1), .CLK(1'b0), .EN(na15_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2905_1_i) );
// C_///AND/D      x115y96     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2906_4 ( .OUT(na2906_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na215_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2906_5 ( .OUT(na2906_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2906_2_i) );
// C_AND/D///      x113y101     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2907_1 ( .OUT(na2907_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na263_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2907_2 ( .OUT(na2907_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2907_1_i) );
// C_///AND/D      x110y73     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2908_4 ( .OUT(na2908_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na275_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2908_5 ( .OUT(na2908_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2908_2_i) );
// C_AND/D///      x112y100     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2909_1 ( .OUT(na2909_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na281_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2909_2 ( .OUT(na2909_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2909_1_i) );
// C_///AND/D      x104y75     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2910_4 ( .OUT(na2910_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na293_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2910_5 ( .OUT(na2910_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2910_2_i) );
// C_AND/D///      x109y81     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2911_1 ( .OUT(na2911_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na298_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2911_2 ( .OUT(na2911_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2911_1_i) );
// C_///AND/D      x107y88     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2912_4 ( .OUT(na2912_2_i), .IN1(na308_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2912_5 ( .OUT(na2912_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2912_2_i) );
// C_AND/D///      x111y82     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2913_1 ( .OUT(na2913_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na312_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2913_2 ( .OUT(na2913_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2913_1_i) );
// C_///AND/D      x131y100     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2914_4 ( .OUT(na2914_2_i), .IN1(na959_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2914_5 ( .OUT(na2914_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2914_2_i) );
// C_AND/D///      x140y101     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2915_1 ( .OUT(na2915_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1003_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2915_2 ( .OUT(na2915_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2915_1_i) );
// C_///AND/D      x136y91     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2916_4 ( .OUT(na2916_2_i), .IN1(na1012_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2916_5 ( .OUT(na2916_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2916_2_i) );
// C_AND/D///      x127y94     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2917_1 ( .OUT(na2917_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1019_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2917_2 ( .OUT(na2917_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2917_1_i) );
// C_///AND/D      x138y79     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2918_4 ( .OUT(na2918_2_i), .IN1(na1025_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2918_5 ( .OUT(na2918_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2918_2_i) );
// C_AND/D///      x126y75     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2919_1 ( .OUT(na2919_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1029_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2919_2 ( .OUT(na2919_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2919_1_i) );
// C_///AND/D      x123y96     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2920_4 ( .OUT(na2920_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1032_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2920_5 ( .OUT(na2920_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2920_2_i) );
// C_AND/D///      x122y81     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2921_1 ( .OUT(na2921_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1034_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2921_2 ( .OUT(na2921_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2921_1_i) );
// C_///AND/D      x138y99     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2922_4 ( .OUT(na2922_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na884_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2922_5 ( .OUT(na2922_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2922_2_i) );
// C_AND/D///      x135y95     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2923_1 ( .OUT(na2923_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na926_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2923_2 ( .OUT(na2923_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2923_1_i) );
// C_///AND/D      x136y82     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2924_4 ( .OUT(na2924_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na935_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2924_5 ( .OUT(na2924_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2924_2_i) );
// C_AND/D///      x137y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2925_1 ( .OUT(na2925_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na941_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2925_2 ( .OUT(na2925_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2925_1_i) );
// C_///AND/D      x132y71     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2926_4 ( .OUT(na2926_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na948_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2926_5 ( .OUT(na2926_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2926_2_i) );
// C_AND/D///      x125y70     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2927_1 ( .OUT(na2927_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na952_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2927_2 ( .OUT(na2927_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2927_1_i) );
// C_///AND/D      x136y80     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2928_4 ( .OUT(na2928_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na955_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2928_5 ( .OUT(na2928_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2928_2_i) );
// C_AND/D///      x130y71     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2929_1 ( .OUT(na2929_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na957_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2929_2 ( .OUT(na2929_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2929_1_i) );
// C_///AND/D      x135y95     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2930_4 ( .OUT(na2930_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na807_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2930_5 ( .OUT(na2930_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2930_2_i) );
// C_///AND/D      x141y96     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2931_4 ( .OUT(na2931_2_i), .IN1(na852_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2931_5 ( .OUT(na2931_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2931_2_i) );
// C_///AND/D      x137y89     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2932_4 ( .OUT(na2932_2_i), .IN1(1'b1), .IN2(na862_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2932_5 ( .OUT(na2932_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2932_2_i) );
// C_AND/D///      x128y93     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2933_1 ( .OUT(na2933_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na866_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2933_2 ( .OUT(na2933_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2933_1_i) );
// C_///AND/D      x137y75     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2934_4 ( .OUT(na2934_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na872_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2934_5 ( .OUT(na2934_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2934_2_i) );
// C_AND/D///      x120y73     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2935_1 ( .OUT(na2935_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na875_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2935_2 ( .OUT(na2935_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2935_1_i) );
// C_///AND/D      x137y86     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2936_4 ( .OUT(na2936_2_i), .IN1(na877_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2936_5 ( .OUT(na2936_2), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2936_2_i) );
// C_AND/D///      x130y77     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2937_1 ( .OUT(na2937_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na881_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2937_2 ( .OUT(na2937_1), .CLK(1'b0), .EN(na1438_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2937_1_i) );
// C_///AND/D      x137y93     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2938_4 ( .OUT(na2938_2_i), .IN1(na1077_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2938_5 ( .OUT(na2938_2), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2938_2_i) );
// C_AND/D///      x137y93     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2939_1 ( .OUT(na2939_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1078_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2939_2 ( .OUT(na2939_1), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2939_1_i) );
// C_///AND/D      x140y84     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2940_4 ( .OUT(na2940_2_i), .IN1(1'b1), .IN2(na1079_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2940_5 ( .OUT(na2940_2), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2940_2_i) );
// C_AND/D///      x133y89     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2941_1 ( .OUT(na2941_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1080_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2941_2 ( .OUT(na2941_1), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2941_1_i) );
// C_///AND/D      x142y77     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2942_4 ( .OUT(na2942_2_i), .IN1(1'b1), .IN2(na1081_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2942_5 ( .OUT(na2942_2), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2942_2_i) );
// C_AND/D///      x133y75     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2943_1 ( .OUT(na2943_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1082_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2943_2 ( .OUT(na2943_1), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2943_1_i) );
// C_///AND/D      x131y89     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2944_4 ( .OUT(na2944_2_i), .IN1(na1083_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2944_5 ( .OUT(na2944_2), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2944_2_i) );
// C_AND/D///      x131y81     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2945_1 ( .OUT(na2945_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1084_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2945_2 ( .OUT(na2945_1), .CLK(1'b0), .EN(na1459_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2945_1_i) );
// C_AND/D//AND/D      x113y74     80'h40_E800_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2946_1 ( .OUT(na2946_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1806_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2946_2 ( .OUT(na2946_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2946_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2946_4 ( .OUT(na2946_2_i), .IN1(na316_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2946_5 ( .OUT(na2946_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2946_2_i) );
// C_AND/D//AND/D      x114y72     80'h40_E800_80_0000_0C88_3FFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2949_1 ( .OUT(na2949_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na285_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2949_2 ( .OUT(na2949_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2949_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2949_4 ( .OUT(na2949_2_i), .IN1(1'b1), .IN2(na354_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2949_5 ( .OUT(na2949_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2949_2_i) );
// C_///AND/D      x112y69     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2950_4 ( .OUT(na2950_2_i), .IN1(1'b1), .IN2(na1821_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2950_5 ( .OUT(na2950_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2950_2_i) );
// C_AND/D//AND/D      x112y71     80'h40_E800_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2953_1 ( .OUT(na2953_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1831_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2953_2 ( .OUT(na2953_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2953_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2953_4 ( .OUT(na2953_2_i), .IN1(na486_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2953_5 ( .OUT(na2953_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2953_2_i) );
// C_AND/D///      x119y73     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2955_1 ( .OUT(na2955_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na327_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2955_2 ( .OUT(na2955_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2955_1_i) );
// C_AND/D//AND/D      x115y74     80'h40_E800_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2956_1 ( .OUT(na2956_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na336_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2956_2 ( .OUT(na2956_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2956_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2956_4 ( .OUT(na2956_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1811_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2956_5 ( .OUT(na2956_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2956_2_i) );
// C_AND/D//AND/D      x113y71     80'h40_E800_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2957_1 ( .OUT(na2957_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na345_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2957_2 ( .OUT(na2957_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2957_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2957_4 ( .OUT(na2957_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na522_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2957_5 ( .OUT(na2957_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2957_2_i) );
// C_AND/D//AND/D      x117y67     80'h40_E800_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2959_1 ( .OUT(na2959_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na363_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2959_2 ( .OUT(na2959_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2959_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2959_4 ( .OUT(na2959_2_i), .IN1(na504_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2959_5 ( .OUT(na2959_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2959_2_i) );
// C_AND/D//AND/D      x115y71     80'h40_E800_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2961_1 ( .OUT(na2961_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na381_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2961_2 ( .OUT(na2961_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2961_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2961_4 ( .OUT(na2961_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1816_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2961_5 ( .OUT(na2961_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2961_2_i) );
// C_///AND/D      x124y65     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2963_4 ( .OUT(na2963_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na398_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2963_5 ( .OUT(na2963_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2963_2_i) );
// C_AND/D///      x120y71     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2964_1 ( .OUT(na2964_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na407_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2964_2 ( .OUT(na2964_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2964_1_i) );
// C_AND/D//AND/D      x117y72     80'h40_E800_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2965_1 ( .OUT(na2965_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na416_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2965_2 ( .OUT(na2965_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2965_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2965_4 ( .OUT(na2965_2_i), .IN1(1'b1), .IN2(na477_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2965_5 ( .OUT(na2965_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2965_2_i) );
// C_AND/D//AND/D      x115y70     80'h40_E800_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2966_1 ( .OUT(na2966_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na425_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2966_2 ( .OUT(na2966_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2966_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2966_4 ( .OUT(na2966_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na495_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2966_5 ( .OUT(na2966_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2966_2_i) );
// C_AND/D//AND/D      x116y67     80'h40_E800_80_0000_0C88_AFF3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2967_1 ( .OUT(na2967_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na434_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2967_2 ( .OUT(na2967_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2967_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2967_4 ( .OUT(na2967_2_i), .IN1(1'b1), .IN2(~na300_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2967_5 ( .OUT(na2967_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2967_2_i) );
// C_AND/D//AND/D      x120y68     80'h40_E800_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2968_1 ( .OUT(na2968_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na442_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2968_2 ( .OUT(na2968_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2968_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2968_4 ( .OUT(na2968_2_i), .IN1(1'b1), .IN2(na372_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2968_5 ( .OUT(na2968_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2968_2_i) );
// C_AND/D//AND/D      x116y72     80'h40_E800_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2969_1 ( .OUT(na2969_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na451_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2969_2 ( .OUT(na2969_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2969_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2969_4 ( .OUT(na2969_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na390_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2969_5 ( .OUT(na2969_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2969_2_i) );
// C_///AND/D      x118y69     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2970_4 ( .OUT(na2970_2_i), .IN1(1'b1), .IN2(na460_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2970_5 ( .OUT(na2970_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2970_2_i) );
// C_AND/D///      x120y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2971_1 ( .OUT(na2971_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na469_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2971_2 ( .OUT(na2971_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2971_1_i) );
// C_AND/D//AND/D      x117y68     80'h40_E800_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2976_1 ( .OUT(na2976_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na513_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2976_2 ( .OUT(na2976_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2976_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2976_4 ( .OUT(na2976_2_i), .IN1(1'b1), .IN2(na1826_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2976_5 ( .OUT(na2976_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2976_2_i) );
// C_///AND/D      x142y91     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2978_4 ( .OUT(na2978_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1037_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2978_5 ( .OUT(na2978_2), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2978_2_i) );
// C_AND/D///      x140y91     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2979_1 ( .OUT(na2979_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1038_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2979_2 ( .OUT(na2979_1), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2979_1_i) );
// C_///AND/D      x141y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2980_4 ( .OUT(na2980_2_i), .IN1(1'b1), .IN2(na1039_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2980_5 ( .OUT(na2980_2), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2980_2_i) );
// C_AND/D///      x138y83     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2981_1 ( .OUT(na2981_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1040_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2981_2 ( .OUT(na2981_1), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2981_1_i) );
// C_///AND/D      x141y74     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2982_4 ( .OUT(na2982_2_i), .IN1(1'b1), .IN2(na1041_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2982_5 ( .OUT(na2982_2), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2982_2_i) );
// C_AND/D///      x138y67     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2983_1 ( .OUT(na2983_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1042_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2983_2 ( .OUT(na2983_1), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2983_1_i) );
// C_///AND/D      x139y79     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2984_4 ( .OUT(na2984_2_i), .IN1(na1043_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2984_5 ( .OUT(na2984_2), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2984_2_i) );
// C_AND/D///      x137y71     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2985_1 ( .OUT(na2985_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1044_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2985_2 ( .OUT(na2985_1), .CLK(1'b0), .EN(na1439_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2985_1_i) );
// C_///AND/D      x142y93     80'h40_E400_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2986_4 ( .OUT(na2986_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1045_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2986_5 ( .OUT(na2986_2), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2986_2_i) );
// C_///AND/D      x141y93     80'h40_E400_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2987_4 ( .OUT(na2987_2_i), .IN1(1'b1), .IN2(na1046_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2987_5 ( .OUT(na2987_2), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2987_2_i) );
// C_///AND/D      x141y71     80'h40_E400_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2988_4 ( .OUT(na2988_2_i), .IN1(1'b1), .IN2(na1047_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2988_5 ( .OUT(na2988_2), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2988_2_i) );
// C_AND/D///      x141y79     80'h40_E400_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2989_1 ( .OUT(na2989_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1048_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2989_2 ( .OUT(na2989_1), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2989_1_i) );
// C_///AND/D      x140y66     80'h40_E400_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2990_4 ( .OUT(na2990_2_i), .IN1(na1049_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2990_5 ( .OUT(na2990_2), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2990_2_i) );
// C_AND/D///      x140y66     80'h40_E400_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2991_1 ( .OUT(na2991_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1050_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2991_2 ( .OUT(na2991_1), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2991_1_i) );
// C_///AND/D      x140y69     80'h40_E400_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2992_4 ( .OUT(na2992_2_i), .IN1(na1051_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2992_5 ( .OUT(na2992_2), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2992_2_i) );
// C_AND/D///      x140y69     80'h40_E400_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2993_1 ( .OUT(na2993_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1052_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2993_2 ( .OUT(na2993_1), .CLK(1'b0), .EN(~na1440_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2993_1_i) );
// C_///AND/D      x137y87     80'h40_E400_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2994_4 ( .OUT(na2994_2_i), .IN1(1'b1), .IN2(na1061_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2994_5 ( .OUT(na2994_2), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2994_2_i) );
// C_AND/D///      x140y92     80'h40_E400_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2995_1 ( .OUT(na2995_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1062_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2995_2 ( .OUT(na2995_1), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2995_1_i) );
// C_///AND/D      x144y80     80'h40_E400_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2996_4 ( .OUT(na2996_2_i), .IN1(na1063_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2996_5 ( .OUT(na2996_2), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2996_2_i) );
// C_AND/D///      x137y87     80'h40_E400_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2997_1 ( .OUT(na2997_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1064_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2997_2 ( .OUT(na2997_1), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2997_1_i) );
// C_///AND/D      x137y73     80'h40_E400_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2998_4 ( .OUT(na2998_2_i), .IN1(1'b1), .IN2(na1065_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2998_5 ( .OUT(na2998_2), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2998_2_i) );
// C_AND/D///      x135y72     80'h40_E400_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2999_1 ( .OUT(na2999_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1066_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2999_2 ( .OUT(na2999_1), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2999_1_i) );
// C_///AND/D      x144y77     80'h40_E400_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3000_4 ( .OUT(na3000_2_i), .IN1(1'b1), .IN2(na1067_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3000_5 ( .OUT(na3000_2), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3000_2_i) );
// C_AND/D///      x134y76     80'h40_E400_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3001_1 ( .OUT(na3001_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1068_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3001_2 ( .OUT(na3001_1), .CLK(1'b0), .EN(~na1442_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3001_1_i) );
// C_///AND/D      x141y92     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3002_4 ( .OUT(na3002_2_i), .IN1(na851_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3002_5 ( .OUT(na3002_2), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3002_2_i) );
// C_AND/D///      x140y88     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3003_1 ( .OUT(na3003_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na861_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3003_2 ( .OUT(na3003_1), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3003_1_i) );
// C_///AND/D      x142y84     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3004_4 ( .OUT(na3004_2_i), .IN1(1'b1), .IN2(na865_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3004_5 ( .OUT(na3004_2), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3004_2_i) );
// C_AND/D///      x139y85     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3005_1 ( .OUT(na3005_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na871_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3005_2 ( .OUT(na3005_1), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3005_1_i) );
// C_///AND/D      x138y68     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3006_4 ( .OUT(na3006_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na874_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3006_5 ( .OUT(na3006_2), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3006_2_i) );
// C_AND/D///      x138y68     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3007_1 ( .OUT(na3007_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na876_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3007_2 ( .OUT(na3007_1), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3007_1_i) );
// C_///AND/D      x143y75     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3008_4 ( .OUT(na3008_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na880_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3008_5 ( .OUT(na3008_2), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3008_2_i) );
// C_AND/D///      x139y70     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3009_1 ( .OUT(na3009_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na883_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3009_2 ( .OUT(na3009_1), .CLK(1'b0), .EN(na1443_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3009_1_i) );
// C_///AND/D      x131y109     80'h40_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3010_4 ( .OUT(na3010_2_i), .IN1(1'b1), .IN2(na1135_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3010_5 ( .OUT(na3010_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3010_2_i) );
// C_AND/D///      x134y109     80'h40_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3011_1 ( .OUT(na3011_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3011_2 ( .OUT(na3011_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3011_1_i) );
// C_///AND/D      x131y110     80'h40_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3013_4 ( .OUT(na3013_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1142_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3013_5 ( .OUT(na3013_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3013_2_i) );
// C_AND/D///      x127y112     80'h40_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3014_1 ( .OUT(na3014_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3014_2 ( .OUT(na3014_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3014_1_i) );
// C_///AND/D      x136y109     80'h40_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3015_4 ( .OUT(na3015_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1146_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3015_5 ( .OUT(na3015_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3015_2_i) );
// C_AND/D///      x131y109     80'h40_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3016_1 ( .OUT(na3016_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1148_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3016_2 ( .OUT(na3016_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3016_1_i) );
// C_AND/D//AND/D      x125y109     80'h40_EC00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3017_1 ( .OUT(na3017_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1150_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3017_2 ( .OUT(na3017_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3017_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3017_4 ( .OUT(na3017_2_i), .IN1(1'b1), .IN2(na1140_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3017_5 ( .OUT(na3017_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3017_2_i) );
// C_AND/D///      x134y105     80'h40_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3018_1 ( .OUT(na3018_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1152_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3018_2 ( .OUT(na3018_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3018_1_i) );
// C_AND/D///      x148y107     80'h40_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3019_1 ( .OUT(na3019_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1154_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3019_2 ( .OUT(na3019_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3019_1_i) );
// C_///AND/D      x138y111     80'h40_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3021_4 ( .OUT(na3021_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1158_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3021_5 ( .OUT(na3021_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3021_2_i) );
// C_AND/D///      x127y96     80'h40_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3022_1 ( .OUT(na3022_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1160_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3022_2 ( .OUT(na3022_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3022_1_i) );
// C_///AND/D      x146y107     80'h40_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3023_4 ( .OUT(na3023_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1162_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3023_5 ( .OUT(na3023_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3023_2_i) );
// C_AND/D///      x139y103     80'h40_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3024_1 ( .OUT(na3024_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1164_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3024_2 ( .OUT(na3024_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3024_1_i) );
// C_AND/D//AND/D      x137y105     80'h40_EC00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3025_1 ( .OUT(na3025_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1166_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3025_2 ( .OUT(na3025_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3025_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3025_4 ( .OUT(na3025_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1156_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3025_5 ( .OUT(na3025_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3025_2_i) );
// C_///AND/D      x146y105     80'h40_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3026_4 ( .OUT(na3026_2_i), .IN1(na1168_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3026_5 ( .OUT(na3026_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3026_2_i) );
// C_AND/D///      x143y101     80'h40_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3027_1 ( .OUT(na3027_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1170_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3027_2 ( .OUT(na3027_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3027_1_i) );
// C_///AND/D      x143y100     80'h40_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3029_4 ( .OUT(na3029_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3029_5 ( .OUT(na3029_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3029_2_i) );
// C_AND/D///      x146y99     80'h40_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3030_1 ( .OUT(na3030_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1176_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3030_2 ( .OUT(na3030_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3030_1_i) );
// C_///AND/D      x138y102     80'h40_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3031_4 ( .OUT(na3031_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1178_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3031_5 ( .OUT(na3031_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3031_2_i) );
// C_AND/D///      x142y100     80'h40_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3032_1 ( .OUT(na3032_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1180_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3032_2 ( .OUT(na3032_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3032_1_i) );
// C_AND/D//AND/D      x140y104     80'h40_EC00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3033_1 ( .OUT(na3033_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1182_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3033_2 ( .OUT(na3033_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3033_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3033_4 ( .OUT(na3033_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1172_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3033_5 ( .OUT(na3033_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3033_2_i) );
// C_///AND/D      x135y113     80'h40_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3034_4 ( .OUT(na3034_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1184_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3034_5 ( .OUT(na3034_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3034_2_i) );
// C_AND/D///      x139y112     80'h40_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3035_1 ( .OUT(na3035_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1186_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3035_2 ( .OUT(na3035_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3035_1_i) );
// C_///AND/D      x140y109     80'h40_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3037_4 ( .OUT(na3037_2_i), .IN1(na1190_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3037_5 ( .OUT(na3037_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3037_2_i) );
// C_AND/D///      x141y112     80'h40_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3038_1 ( .OUT(na3038_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1192_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3038_2 ( .OUT(na3038_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3038_1_i) );
// C_///AND/D      x139y111     80'h40_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3039_4 ( .OUT(na3039_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1194_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3039_5 ( .OUT(na3039_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3039_2_i) );
// C_AND/D///      x141y111     80'h40_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3040_1 ( .OUT(na3040_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1196_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3040_2 ( .OUT(na3040_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3040_1_i) );
// C_AND/D//AND/D      x138y112     80'h40_EC00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3041_1 ( .OUT(na3041_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1198_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3041_2 ( .OUT(na3041_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3041_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3041_4 ( .OUT(na3041_2_i), .IN1(na1188_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3041_5 ( .OUT(na3041_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3041_2_i) );
// C_///AND/D      x139y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3042_4 ( .OUT(na3042_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na925_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3042_5 ( .OUT(na3042_2), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3042_2_i) );
// C_AND/D///      x138y85     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3043_1 ( .OUT(na3043_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na934_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3043_2 ( .OUT(na3043_1), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3043_1_i) );
// C_///AND/D      x144y74     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3044_4 ( .OUT(na3044_2_i), .IN1(na940_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3044_5 ( .OUT(na3044_2), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3044_2_i) );
// C_AND/D///      x141y87     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3045_1 ( .OUT(na3045_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na947_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3045_2 ( .OUT(na3045_1), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3045_1_i) );
// C_///AND/D      x139y68     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3046_4 ( .OUT(na3046_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na951_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3046_5 ( .OUT(na3046_2), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3046_2_i) );
// C_AND/D///      x140y67     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3047_1 ( .OUT(na3047_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na954_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3047_2 ( .OUT(na3047_1), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3047_1_i) );
// C_///AND/D      x139y75     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3048_4 ( .OUT(na3048_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na956_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3048_5 ( .OUT(na3048_2), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3048_2_i) );
// C_AND/D///      x139y68     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3049_1 ( .OUT(na3049_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na958_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3049_2 ( .OUT(na3049_1), .CLK(1'b0), .EN(na1447_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3049_1_i) );
// C_///AND/D      x138y91     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3050_4 ( .OUT(na3050_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1053_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3050_5 ( .OUT(na3050_2), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3050_2_i) );
// C_AND/D///      x139y91     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3051_1 ( .OUT(na3051_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1054_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3051_2 ( .OUT(na3051_1), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3051_1_i) );
// C_///AND/D      x139y81     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3052_4 ( .OUT(na3052_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1055_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3052_5 ( .OUT(na3052_2), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3052_2_i) );
// C_AND/D///      x133y85     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3053_1 ( .OUT(na3053_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1056_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3053_2 ( .OUT(na3053_1), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3053_1_i) );
// C_AND/D///      x140y75     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3054_1 ( .OUT(na3054_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1057_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3054_2 ( .OUT(na3054_1), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3054_1_i) );
// C_AND/D///      x138y69     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3055_1 ( .OUT(na3055_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1058_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3055_2 ( .OUT(na3055_1), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3055_1_i) );
// C_///AND/D      x140y81     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3056_4 ( .OUT(na3056_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1059_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3056_5 ( .OUT(na3056_2), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3056_2_i) );
// C_AND/D///      x133y77     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3057_1 ( .OUT(na3057_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1060_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3057_2 ( .OUT(na3057_1), .CLK(1'b0), .EN(na1445_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3057_1_i) );
// C_///AND/D      x140y89     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3058_4 ( .OUT(na3058_2_i), .IN1(1'b1), .IN2(na1002_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3058_5 ( .OUT(na3058_2), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3058_2_i) );
// C_AND/D///      x140y90     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3059_1 ( .OUT(na3059_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1011_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3059_2 ( .OUT(na3059_1), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3059_1_i) );
// C_///AND/D      x138y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3060_4 ( .OUT(na3060_2_i), .IN1(1'b1), .IN2(na1018_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3060_5 ( .OUT(na3060_2), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3060_2_i) );
// C_AND/D///      x135y91     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3061_1 ( .OUT(na3061_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1024_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3061_2 ( .OUT(na3061_1), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3061_1_i) );
// C_///AND/D      x139y71     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3062_4 ( .OUT(na3062_2_i), .IN1(na1028_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3062_5 ( .OUT(na3062_2), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3062_2_i) );
// C_AND/D///      x139y71     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3063_1 ( .OUT(na3063_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1031_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3063_2 ( .OUT(na3063_1), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3063_1_i) );
// C_///AND/D      x141y84     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3064_4 ( .OUT(na3064_2_i), .IN1(na1033_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3064_5 ( .OUT(na3064_2), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3064_2_i) );
// C_AND/D///      x129y82     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3065_1 ( .OUT(na3065_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1036_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3065_2 ( .OUT(na3065_1), .CLK(1'b0), .EN(na1450_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3065_1_i) );
// C_///AND/D      x138y92     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3066_4 ( .OUT(na3066_2_i), .IN1(1'b1), .IN2(na1069_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3066_5 ( .OUT(na3066_2), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3066_2_i) );
// C_AND/D///      x135y88     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3067_1 ( .OUT(na3067_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1070_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3067_2 ( .OUT(na3067_1), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3067_1_i) );
// C_///AND/D      x140y79     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3068_4 ( .OUT(na3068_2_i), .IN1(na1071_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3068_5 ( .OUT(na3068_2), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3068_2_i) );
// C_AND/D///      x137y90     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3069_1 ( .OUT(na3069_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1072_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3069_2 ( .OUT(na3069_1), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3069_1_i) );
// C_///AND/D      x139y67     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3070_4 ( .OUT(na3070_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1073_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3070_5 ( .OUT(na3070_2), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3070_2_i) );
// C_AND/D///      x134y70     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3071_1 ( .OUT(na3071_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1074_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3071_2 ( .OUT(na3071_1), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3071_1_i) );
// C_///AND/D      x133y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3072_4 ( .OUT(na3072_2_i), .IN1(1'b1), .IN2(na1075_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3072_5 ( .OUT(na3072_2), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3072_2_i) );
// C_AND/D///      x134y74     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3073_1 ( .OUT(na3073_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1076_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3073_2 ( .OUT(na3073_1), .CLK(1'b0), .EN(na1446_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3073_1_i) );
// C_///AND/D      x139y93     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3074_4 ( .OUT(na3074_2_i), .IN1(na1109_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3074_5 ( .OUT(na3074_2), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3074_2_i) );
// C_AND/D///      x137y92     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3075_1 ( .OUT(na3075_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1110_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3075_2 ( .OUT(na3075_1), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3075_1_i) );
// C_///AND/D      x141y85     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3076_4 ( .OUT(na3076_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1111_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3076_5 ( .OUT(na3076_2), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3076_2_i) );
// C_AND/D///      x134y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3077_1 ( .OUT(na3077_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1112_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3077_2 ( .OUT(na3077_1), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3077_1_i) );
// C_///AND/D      x143y77     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3078_4 ( .OUT(na3078_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1113_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3078_5 ( .OUT(na3078_2), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3078_2_i) );
// C_AND/D///      x134y72     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3079_1 ( .OUT(na3079_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1114_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3079_2 ( .OUT(na3079_1), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3079_1_i) );
// C_///AND/D      x138y86     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3080_4 ( .OUT(na3080_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1115_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3080_5 ( .OUT(na3080_2), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3080_2_i) );
// C_AND/D///      x132y78     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3081_1 ( .OUT(na3081_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1116_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3081_2 ( .OUT(na3081_1), .CLK(1'b0), .EN(na1452_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3081_1_i) );
// C_///AND/D      x141y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3082_4 ( .OUT(na3082_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1101_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3082_5 ( .OUT(na3082_2), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3082_2_i) );
// C_///AND/D      x138y89     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3083_4 ( .OUT(na3083_2_i), .IN1(1'b1), .IN2(na1102_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3083_5 ( .OUT(na3083_2), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3083_2_i) );
// C_///AND/D      x138y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3084_4 ( .OUT(na3084_2_i), .IN1(1'b1), .IN2(na1103_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3084_5 ( .OUT(na3084_2), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3084_2_i) );
// C_AND/D///      x140y87     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3085_1 ( .OUT(na3085_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1104_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3085_2 ( .OUT(na3085_1), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3085_1_i) );
// C_///AND/D      x141y69     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3086_4 ( .OUT(na3086_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1105_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3086_5 ( .OUT(na3086_2), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3086_2_i) );
// C_AND/D///      x137y67     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3087_1 ( .OUT(na3087_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1106_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3087_2 ( .OUT(na3087_1), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3087_1_i) );
// C_///AND/D      x139y69     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3088_4 ( .OUT(na3088_2_i), .IN1(na1107_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3088_5 ( .OUT(na3088_2), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3088_2_i) );
// C_AND/D///      x137y69     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3089_1 ( .OUT(na3089_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1108_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3089_2 ( .OUT(na3089_1), .CLK(1'b0), .EN(na1449_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3089_1_i) );
// C_///AND/D      x132y87     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3090_4 ( .OUT(na3090_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1085_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3090_5 ( .OUT(na3090_2), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3090_2_i) );
// C_AND/D///      x136y93     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3091_1 ( .OUT(na3091_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1086_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3091_2 ( .OUT(na3091_1), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3091_1_i) );
// C_///AND/D      x136y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3092_4 ( .OUT(na3092_2_i), .IN1(1'b1), .IN2(na1087_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3092_5 ( .OUT(na3092_2), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3092_2_i) );
// C_AND/D///      x132y87     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3093_1 ( .OUT(na3093_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1088_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3093_2 ( .OUT(na3093_1), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3093_1_i) );
// C_///AND/D      x135y74     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3094_4 ( .OUT(na3094_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1089_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3094_5 ( .OUT(na3094_2), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3094_2_i) );
// C_AND/D///      x135y78     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3095_1 ( .OUT(na3095_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1090_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3095_2 ( .OUT(na3095_1), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3095_1_i) );
// C_///AND/D      x134y81     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3096_4 ( .OUT(na3096_2_i), .IN1(na1091_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3096_5 ( .OUT(na3096_2), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3096_2_i) );
// C_AND/D///      x135y77     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3097_1 ( .OUT(na3097_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1092_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3097_2 ( .OUT(na3097_1), .CLK(1'b0), .EN(na1451_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3097_1_i) );
// C_///AND/D      x114y92     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3098_4 ( .OUT(na3098_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na13_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3098_5 ( .OUT(na3098_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3098_2_i) );
// C_AND/D///      x121y94     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3099_1 ( .OUT(na3099_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na28_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3099_2 ( .OUT(na3099_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3099_1_i) );
// C_///AND/D      x116y77     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3100_4 ( .OUT(na3100_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na34_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3100_5 ( .OUT(na3100_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3100_2_i) );
// C_AND/D///      x107y98     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3101_1 ( .OUT(na3101_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na40_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3101_2 ( .OUT(na3101_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3101_1_i) );
// C_///AND/D      x106y72     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3102_4 ( .OUT(na3102_2_i), .IN1(na46_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3102_5 ( .OUT(na3102_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3102_2_i) );
// C_AND/D///      x112y75     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3103_1 ( .OUT(na3103_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na52_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3103_2 ( .OUT(na3103_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3103_1_i) );
// C_///AND/D      x108y80     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3104_4 ( .OUT(na3104_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na59_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3104_5 ( .OUT(na3104_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3104_2_i) );
// C_AND/D///      x108y68     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3105_1 ( .OUT(na3105_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na65_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3105_2 ( .OUT(na3105_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3105_1_i) );
// C_///AND/D      x134y97     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3106_4 ( .OUT(na3106_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na71_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3106_5 ( .OUT(na3106_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3106_2_i) );
// C_AND/D///      x139y96     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3107_1 ( .OUT(na3107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na77_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3107_2 ( .OUT(na3107_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3107_1_i) );
// C_///AND/D      x133y91     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3108_4 ( .OUT(na3108_2_i), .IN1(na83_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3108_5 ( .OUT(na3108_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3108_2_i) );
// C_AND/D///      x124y96     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3109_1 ( .OUT(na3109_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na89_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3109_2 ( .OUT(na3109_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3109_1_i) );
// C_///AND/D      x136y77     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3110_4 ( .OUT(na3110_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na95_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3110_5 ( .OUT(na3110_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3110_2_i) );
// C_AND/D///      x120y78     80'h40_E800_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3111_1 ( .OUT(na3111_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na101_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3111_2 ( .OUT(na3111_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3111_1_i) );
// C_///AND/D      x131y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3112_4 ( .OUT(na3112_2_i), .IN1(1'b1), .IN2(na107_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3112_5 ( .OUT(na3112_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3112_2_i) );
// C_///AND/D      x112y73     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3113_4 ( .OUT(na3113_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na113_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3113_5 ( .OUT(na3113_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3113_2_i) );
// C_///AND/D      x133y95     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3114_4 ( .OUT(na3114_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na119_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3114_5 ( .OUT(na3114_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3114_2_i) );
// C_AND/D///      x140y93     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3115_1 ( .OUT(na3115_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na125_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3115_2 ( .OUT(na3115_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3115_1_i) );
// C_///AND/D      x134y89     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3116_4 ( .OUT(na3116_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na131_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3116_5 ( .OUT(na3116_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3116_2_i) );
// C_AND/D///      x128y96     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3117_1 ( .OUT(na3117_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na137_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3117_2 ( .OUT(na3117_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3117_1_i) );
// C_///AND/D      x128y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3118_4 ( .OUT(na3118_2_i), .IN1(1'b1), .IN2(na143_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3118_5 ( .OUT(na3118_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3118_2_i) );
// C_AND/D///      x117y73     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3119_1 ( .OUT(na3119_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na149_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3119_2 ( .OUT(na3119_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3119_1_i) );
// C_///AND/D      x130y75     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3120_4 ( .OUT(na3120_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na155_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3120_5 ( .OUT(na3120_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3120_2_i) );
// C_AND/D///      x118y78     80'h40_E800_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3121_1 ( .OUT(na3121_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na161_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3121_2 ( .OUT(na3121_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3121_1_i) );
// C_///AND/D      x123y104     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3122_4 ( .OUT(na3122_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na167_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3122_5 ( .OUT(na3122_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3122_2_i) );
// C_AND/D///      x133y98     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3123_1 ( .OUT(na3123_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na173_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3123_2 ( .OUT(na3123_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3123_1_i) );
// C_///AND/D      x128y95     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3124_4 ( .OUT(na3124_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na179_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3124_5 ( .OUT(na3124_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3124_2_i) );
// C_AND/D///      x118y96     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3125_1 ( .OUT(na3125_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na185_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3125_2 ( .OUT(na3125_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3125_1_i) );
// C_///AND/D      x121y83     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3126_4 ( .OUT(na3126_2_i), .IN1(1'b1), .IN2(na191_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3126_5 ( .OUT(na3126_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3126_2_i) );
// C_AND/D///      x116y82     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3127_1 ( .OUT(na3127_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na197_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3127_2 ( .OUT(na3127_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3127_1_i) );
// C_///AND/D      x118y89     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3128_4 ( .OUT(na3128_2_i), .IN1(1'b1), .IN2(na203_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3128_5 ( .OUT(na3128_2), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3128_2_i) );
// C_AND/D///      x111y86     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3129_1 ( .OUT(na3129_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na209_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3129_2 ( .OUT(na3129_1), .CLK(1'b0), .EN(na543_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3129_1_i) );
// C_///AND/D      x122y73     80'h40_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3130_4 ( .OUT(na3130_2_i), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3130_5 ( .OUT(na3130_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3130_2_i) );
// C_AND/D///      x127y65     80'h40_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3131_1 ( .OUT(na3131_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2415_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3131_2 ( .OUT(na3131_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3131_1_i) );
// C_///AND/D      x125y74     80'h40_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3132_4 ( .OUT(na3132_2_i), .IN1(1'b1), .IN2(na2416_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3132_5 ( .OUT(na3132_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3132_2_i) );
// C_AND/D///      x125y66     80'h40_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3133_1 ( .OUT(na3133_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2417_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3133_2 ( .OUT(na3133_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3133_1_i) );
// C_///AND/D      x134y83     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3134_4 ( .OUT(na3134_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1117_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3134_5 ( .OUT(na3134_2), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3134_2_i) );
// C_AND/D///      x130y86     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3135_1 ( .OUT(na3135_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1118_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3135_2 ( .OUT(na3135_1), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3135_1_i) );
// C_///AND/D      x131y76     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3136_4 ( .OUT(na3136_2_i), .IN1(na1119_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3136_5 ( .OUT(na3136_2), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3136_2_i) );
// C_AND/D///      x126y85     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3137_1 ( .OUT(na3137_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1120_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3137_2 ( .OUT(na3137_1), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3137_1_i) );
// C_///AND/D      x128y72     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3138_4 ( .OUT(na3138_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1121_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3138_5 ( .OUT(na3138_2), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3138_2_i) );
// C_AND/D///      x127y70     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3139_1 ( .OUT(na3139_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1122_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3139_2 ( .OUT(na3139_1), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3139_1_i) );
// C_///AND/D      x127y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3140_4 ( .OUT(na3140_2_i), .IN1(1'b1), .IN2(na1123_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3140_5 ( .OUT(na3140_2), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3140_2_i) );
// C_AND/D///      x127y69     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3141_1 ( .OUT(na3141_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1124_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3141_2 ( .OUT(na3141_1), .CLK(1'b0), .EN(na1458_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3141_1_i) );
// C_AND/D///      x91y105     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3142_1 ( .OUT(na3142_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3142_2 ( .OUT(na3142_1), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3142_1_i) );
// C_AND/D///      x117y111     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3143_1 ( .OUT(na3143_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3143_2 ( .OUT(na3143_1), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3143_1_i) );
// C_///AND/D      x101y93     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3144_4 ( .OUT(na3144_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3144_5 ( .OUT(na3144_2), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3144_2_i) );
// C_AND/D///      x94y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3145_1 ( .OUT(na3145_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3145_2 ( .OUT(na3145_1), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3145_1_i) );
// C_///AND/D      x91y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3146_4 ( .OUT(na3146_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3146_5 ( .OUT(na3146_2), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3146_2_i) );
// C_AND/D///      x94y76     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3147_1 ( .OUT(na3147_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3147_2 ( .OUT(na3147_1), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3147_1_i) );
// C_///AND/D      x91y90     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3148_4 ( .OUT(na3148_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3148_5 ( .OUT(na3148_2), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3148_2_i) );
// C_AND/D///      x93y66     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3149_1 ( .OUT(na3149_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3149_2 ( .OUT(na3149_1), .CLK(1'b0), .EN(na1466_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3149_1_i) );
// C_///AND/D      x126y72     80'h40_EC00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3150_4 ( .OUT(na3150_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1317_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3150_5 ( .OUT(na3150_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3150_2_i) );
// C_AND/DST//AND/DST      x126y71     80'h60_BC00_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3151_1 ( .OUT(na3151_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1318_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0100)) 
           _a3151_2 ( .OUT(na3151_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3151_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3151_4 ( .OUT(na3151_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1850_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0100)) 
           _a3151_5 ( .OUT(na3151_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3151_2_i) );
// C_AND/D///      x87y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3153_1 ( .OUT(na3153_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3153_2 ( .OUT(na3153_1), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3153_1_i) );
// C_///AND/D      x118y113     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3154_4 ( .OUT(na3154_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3154_5 ( .OUT(na3154_2), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3154_2_i) );
// C_AND/D///      x102y96     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3155_1 ( .OUT(na3155_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3155_2 ( .OUT(na3155_1), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3155_1_i) );
// C_///AND/D      x88y114     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3156_4 ( .OUT(na3156_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3156_5 ( .OUT(na3156_2), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3156_2_i) );
// C_AND/D///      x91y91     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3157_1 ( .OUT(na3157_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3157_2 ( .OUT(na3157_1), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3157_1_i) );
// C_///AND/D      x91y68     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3158_4 ( .OUT(na3158_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3158_5 ( .OUT(na3158_2), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3158_2_i) );
// C_AND/D///      x91y89     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3159_1 ( .OUT(na3159_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3159_2 ( .OUT(na3159_1), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3159_1_i) );
// C_///AND/D      x92y65     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3160_4 ( .OUT(na3160_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3160_5 ( .OUT(na3160_2), .CLK(1'b0), .EN(na1464_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3160_2_i) );
// C_AND/D///      x98y105     80'h40_F800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3161_1 ( .OUT(na3161_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3161_2 ( .OUT(na3161_1), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3161_1_i) );
// C_///AND/D      x116y105     80'h40_F800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3162_4 ( .OUT(na3162_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3162_5 ( .OUT(na3162_2), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3162_2_i) );
// C_AND/D///      x102y102     80'h40_F800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3163_1 ( .OUT(na3163_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3163_2 ( .OUT(na3163_1), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3163_1_i) );
// C_///AND/D      x98y110     80'h40_F800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3164_4 ( .OUT(na3164_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3164_5 ( .OUT(na3164_2), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3164_2_i) );
// C_AND/D///      x100y92     80'h40_F800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3165_1 ( .OUT(na3165_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3165_2 ( .OUT(na3165_1), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3165_1_i) );
// C_///AND/D      x102y71     80'h40_F800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3166_4 ( .OUT(na3166_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3166_5 ( .OUT(na3166_2), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3166_2_i) );
// C_AND/D///      x93y90     80'h40_F800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3167_1 ( .OUT(na3167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3167_2 ( .OUT(na3167_1), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3167_1_i) );
// C_///AND/D      x93y71     80'h40_F800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3168_4 ( .OUT(na3168_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3211_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3168_5 ( .OUT(na3168_2), .CLK(1'b0), .EN(na1381_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3168_2_i) );
// C_AND/D///      x90y103     80'h40_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3169_1 ( .OUT(na3169_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1323_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3169_2 ( .OUT(na3169_1), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3169_1_i) );
// C_AND/D//AND/D      x90y67     80'h40_E800_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3170_1 ( .OUT(na3170_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1329_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3170_2 ( .OUT(na3170_1), .CLK(1'b0), .EN(na1435_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3170_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3170_4 ( .OUT(na3170_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1330_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3170_5 ( .OUT(na3170_2), .CLK(1'b0), .EN(na1435_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3170_2_i) );
// C_///AND/D      x90y68     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3172_4 ( .OUT(na3172_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1331_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3172_5 ( .OUT(na3172_2), .CLK(1'b0), .EN(na1435_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3172_2_i) );
// C_AND/D///      x88y68     80'h40_E400_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3173_1 ( .OUT(na3173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1332_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3173_2 ( .OUT(na3173_1), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3173_1_i) );
// C_///AND/D      x90y69     80'h40_E400_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3174_4 ( .OUT(na3174_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1337_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3174_5 ( .OUT(na3174_2), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3174_2_i) );
// C_AND/D//AND/D      x89y67     80'h40_E400_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3175_1 ( .OUT(na3175_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1338_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3175_2 ( .OUT(na3175_1), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3175_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3175_4 ( .OUT(na3175_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1340_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3175_5 ( .OUT(na3175_2), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3175_2_i) );
// C_AND/D///      x87y68     80'h40_E400_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3176_1 ( .OUT(na3176_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1339_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3176_2 ( .OUT(na3176_1), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3176_1_i) );
// C_AND/D///      x87y69     80'h40_E400_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3178_1 ( .OUT(na3178_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3178_2 ( .OUT(na3178_1), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3178_1_i) );
// C_AND/D///      x88y71     80'h40_E400_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3180_1 ( .OUT(na3180_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1343_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3180_2 ( .OUT(na3180_1), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3180_1_i) );
// C_AND/D//AND/D      x87y76     80'h40_E400_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3181_1 ( .OUT(na3181_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1344_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3181_2 ( .OUT(na3181_1), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3181_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3181_4 ( .OUT(na3181_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1346_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3181_5 ( .OUT(na3181_2), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3181_2_i) );
// C_AND/D//AND/D      x90y72     80'h40_E400_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3182_1 ( .OUT(na3182_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1345_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3182_2 ( .OUT(na3182_1), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3182_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3182_4 ( .OUT(na3182_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1342_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3182_5 ( .OUT(na3182_2), .CLK(1'b0), .EN(~na1436_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3182_2_i) );
// C_///AND/D      x90y73     80'h40_E800_80_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3184_4 ( .OUT(na3184_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3184_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3184_5 ( .OUT(na3184_2), .CLK(1'b0), .EN(na1384_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3184_2_i) );
// C_AND/D///      x89y78     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3185_1 ( .OUT(na3185_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1347_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3185_2 ( .OUT(na3185_1), .CLK(1'b0), .EN(na1384_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3185_1_i) );
// C_///AND/D      x112y110     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3186_4 ( .OUT(na3186_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3186_5 ( .OUT(na3186_2), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3186_2_i) );
// C_AND/D///      x116y100     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3187_1 ( .OUT(na3187_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3187_2 ( .OUT(na3187_1), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3187_1_i) );
// C_///AND/D      x110y96     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3188_4 ( .OUT(na3188_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3188_5 ( .OUT(na3188_2), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3188_2_i) );
// C_AND/D///      x97y100     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3189_1 ( .OUT(na3189_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3189_2 ( .OUT(na3189_1), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3189_1_i) );
// C_///AND/D      x102y86     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3190_4 ( .OUT(na3190_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3190_5 ( .OUT(na3190_2), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3190_2_i) );
// C_AND/D///      x102y74     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3191_1 ( .OUT(na3191_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3191_2 ( .OUT(na3191_1), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3191_1_i) );
// C_///AND/D      x104y84     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3192_4 ( .OUT(na3192_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3192_5 ( .OUT(na3192_2), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3192_2_i) );
// C_AND/D///      x102y80     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3193_1 ( .OUT(na3193_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3193_2 ( .OUT(na3193_1), .CLK(1'b0), .EN(na1386_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3193_1_i) );
// C_///AND/D      x99y109     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3194_4 ( .OUT(na3194_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3161_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3194_5 ( .OUT(na3194_2), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3194_2_i) );
// C_AND/D///      x121y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3195_1 ( .OUT(na3195_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3195_2 ( .OUT(na3195_1), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3195_1_i) );
// C_///AND/D      x111y107     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3196_4 ( .OUT(na3196_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3163_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3196_5 ( .OUT(na3196_2), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3196_2_i) );
// C_AND/D///      x100y108     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3197_1 ( .OUT(na3197_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3164_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3197_2 ( .OUT(na3197_1), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3197_1_i) );
// C_///AND/D      x99y91     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3198_4 ( .OUT(na3198_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3198_5 ( .OUT(na3198_2), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3198_2_i) );
// C_AND/D///      x97y84     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3199_1 ( .OUT(na3199_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3166_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3199_2 ( .OUT(na3199_1), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3199_1_i) );
// C_///AND/D      x99y93     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3200_4 ( .OUT(na3200_2_i), .IN1(1'b1), .IN2(na3167_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3200_5 ( .OUT(na3200_2), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3200_2_i) );
// C_AND/D///      x92y84     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3201_1 ( .OUT(na3201_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3168_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3201_2 ( .OUT(na3201_1), .CLK(1'b0), .EN(na1465_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3201_1_i) );
// C_///AND/D      x99y116     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3202_4 ( .OUT(na3202_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na800_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3202_5 ( .OUT(na3202_2), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3202_2_i) );
// C_AND/D///      x116y115     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3203_1 ( .OUT(na3203_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na799_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3203_2 ( .OUT(na3203_1), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3203_1_i) );
// C_///AND/D      x105y116     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3204_4 ( .OUT(na3204_2_i), .IN1(1'b1), .IN2(na801_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3204_5 ( .OUT(na3204_2), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3204_2_i) );
// C_AND/D///      x99y116     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3205_1 ( .OUT(na3205_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na802_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3205_2 ( .OUT(na3205_1), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3205_1_i) );
// C_///AND/D      x96y116     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3206_4 ( .OUT(na3206_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na803_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3206_5 ( .OUT(na3206_2), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3206_2_i) );
// C_AND/D///      x93y115     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3207_1 ( .OUT(na3207_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na804_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3207_2 ( .OUT(na3207_1), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3207_1_i) );
// C_///AND/D      x87y111     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3208_4 ( .OUT(na3208_2_i), .IN1(na805_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3208_5 ( .OUT(na3208_2), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3208_2_i) );
// C_AND/D///      x90y109     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3209_1 ( .OUT(na3209_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na806_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3209_2 ( .OUT(na3209_1), .CLK(1'b0), .EN(na1441_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3209_1_i) );
// C_///AND/DST      x147y72     80'h60_BC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3210_4 ( .OUT(na3210_2_i), .IN1(na1348_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0100)) 
           _a3210_5 ( .OUT(na3210_2), .CLK(1'b0), .EN(1'b1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3210_2_i) );
// C_///AND/D      x88y76     80'h40_F800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3211_4 ( .OUT(na3211_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3269_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3211_5 ( .OUT(na3211_2), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3211_2_i) );
// C_///AND/D      x146y71     80'h40_F800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3212_4 ( .OUT(na3212_2_i), .IN1(na1356_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3212_5 ( .OUT(na3212_2), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3212_2_i) );
// C_AND/D///      x143y66     80'h40_F800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3213_1 ( .OUT(na3213_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1362_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3213_2 ( .OUT(na3213_1), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3213_1_i) );
// C_AND/D//AND/D      x143y67     80'h40_F800_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3214_1 ( .OUT(na3214_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1363_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3214_2 ( .OUT(na3214_1), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3214_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3214_4 ( .OUT(na3214_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1367_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3214_5 ( .OUT(na3214_2), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3214_2_i) );
// C_///AND/D      x141y67     80'h40_F800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3215_4 ( .OUT(na3215_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1364_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3215_5 ( .OUT(na3215_2), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3215_2_i) );
// C_AND/D//AND/D      x146y69     80'h40_F800_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3216_1 ( .OUT(na3216_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1365_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3216_2 ( .OUT(na3216_1), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3216_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3216_4 ( .OUT(na3216_2_i), .IN1(1'b1), .IN2(na1371_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3216_5 ( .OUT(na3216_2), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3216_2_i) );
// C_AND/D///      x141y68     80'h40_F800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3217_1 ( .OUT(na3217_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1366_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3217_2 ( .OUT(na3217_1), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3217_1_i) );
// C_///AND/D      x142y68     80'h40_F800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3219_4 ( .OUT(na3219_2_i), .IN1(na1368_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3219_5 ( .OUT(na3219_2), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3219_2_i) );
// C_AND/D//AND/D      x144y72     80'h40_F800_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3220_1 ( .OUT(na3220_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1369_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3220_2 ( .OUT(na3220_1), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3220_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3220_4 ( .OUT(na3220_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1370_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3220_5 ( .OUT(na3220_2), .CLK(1'b0), .EN(na3277_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3220_2_i) );
// C_AND/D//AND/D      x148y67     80'h40_E800_80_0000_0C88_5FFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3223_1 ( .OUT(na3223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3223_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3223_2 ( .OUT(na3223_1), .CLK(1'b0), .EN(na1378_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3223_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3223_4 ( .OUT(na3223_2_i), .IN1(1'b1), .IN2(na1372_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3223_5 ( .OUT(na3223_2), .CLK(1'b0), .EN(na1378_1), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3223_2_i) );
// C_AND/D///      x97y107     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3225_1 ( .OUT(na3225_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3161_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3225_2 ( .OUT(na3225_1), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3225_1_i) );
// C_///AND/D      x122y105     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3226_4 ( .OUT(na3226_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3226_5 ( .OUT(na3226_2), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3226_2_i) );
// C_AND/D///      x105y103     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3227_1 ( .OUT(na3227_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3227_2 ( .OUT(na3227_1), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3227_1_i) );
// C_///AND/D      x104y108     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3228_4 ( .OUT(na3228_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3164_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3228_5 ( .OUT(na3228_2), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3228_2_i) );
// C_AND/D///      x101y96     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3229_1 ( .OUT(na3229_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3229_2 ( .OUT(na3229_1), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3229_1_i) );
// C_///AND/D      x97y80     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3230_4 ( .OUT(na3230_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3166_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3230_5 ( .OUT(na3230_2), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3230_2_i) );
// C_AND/D///      x99y96     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3231_1 ( .OUT(na3231_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3167_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3231_2 ( .OUT(na3231_1), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3231_1_i) );
// C_///AND/D      x98y79     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3232_4 ( .OUT(na3232_2_i), .IN1(na3168_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3232_5 ( .OUT(na3232_2), .CLK(1'b0), .EN(na1461_2), .SR(na3277_1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3232_2_i) );
// C_AND/D///      x145y70     80'h40_F800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3234_1 ( .OUT(na3234_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1200_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3234_2 ( .OUT(na3234_1), .CLK(1'b0), .EN(na1383_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3234_1_i) );
// C_AND/D//AND/D      x147y71     80'h40_F800_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3235_1 ( .OUT(na3235_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1201_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3235_2 ( .OUT(na3235_1), .CLK(1'b0), .EN(na1383_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3235_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3235_4 ( .OUT(na3235_2_i), .IN1(1'b1), .IN2(na1202_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3235_5 ( .OUT(na3235_2), .CLK(1'b0), .EN(na1383_1), .SR(1'b1), .CINY2(na4481_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3235_2_i) );
// C_MX2b////      x118y75     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3236_1 ( .OUT(na3236_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1728_1), .IN6(na2946_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y76     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3237_1 ( .OUT(na3237_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1730_1), .IN6(na2956_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y74     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3238_1 ( .OUT(na3238_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2961_2), .IN6(na1733_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y76     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3239_1 ( .OUT(na3239_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1735_1), .IN8(na2949_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y72     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3240_1 ( .OUT(na3240_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2950_2), .IN8(na1737_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y74     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3241_1 ( .OUT(na3241_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2967_2), .IN8(na1739_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y74     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3242_1 ( .OUT(na3242_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1741_1), .IN6(na2976_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y73     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3243_1 ( .OUT(na3243_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2953_1), .IN8(na1743_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y71     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3244_1 ( .OUT(na3244_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1745_2), .IN6(na2946_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y70     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3245_1 ( .OUT(na3245_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4279_2), .IN5(na2955_1), .IN6(1'b0), .IN7(na1746_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y70     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3246_1 ( .OUT(na3246_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1748_1), .IN6(na2956_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y77     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3247_1 ( .OUT(na3247_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2957_1), .IN6(na1750_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y67     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3248_1 ( .OUT(na3248_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1752_1), .IN8(na2949_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y71     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3249_1 ( .OUT(na3249_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2959_1), .IN6(na1754_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y68     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3250_1 ( .OUT(na3250_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1756_1), .IN8(na2968_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3251_1 ( .OUT(na3251_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2961_1), .IN6(na1758_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y70     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3252_1 ( .OUT(na3252_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1760_2), .IN8(na2969_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y68     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3253_1 ( .OUT(na3253_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2963_2), .IN8(na1761_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y69     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3254_1 ( .OUT(na3254_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4279_2), .IN5(na1763_1), .IN6(1'b0), .IN7(na2964_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y70     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3255_1 ( .OUT(na3255_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4279_2), .IN5(1'b0), .IN6(na2965_1), .IN7(1'b0), .IN8(na1765_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y68     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3256_1 ( .OUT(na3256_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4279_2), .IN5(1'b0), .IN6(na2966_1), .IN7(1'b0), .IN8(na1767_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y66     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3257_1 ( .OUT(na3257_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4279_2), .IN5(na1769_1), .IN6(1'b0), .IN7(na2967_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y68     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3258_1 ( .OUT(na3258_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4279_2), .IN5(1'b0), .IN6(na1770_1), .IN7(1'b0), .IN8(na2968_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y65     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3259_1 ( .OUT(na3259_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1771_1), .IN8(na2969_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y72     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3260_1 ( .OUT(na3260_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2970_2), .IN8(na1773_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y69     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3261_1 ( .OUT(na3261_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4279_2), .IN5(1'b0), .IN6(na1775_1), .IN7(1'b0), .IN8(na2971_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y72     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3262_1 ( .OUT(na3262_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1776_2), .IN6(na2965_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y76     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3263_1 ( .OUT(na3263_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2953_2), .IN8(na1777_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y70     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3264_1 ( .OUT(na3264_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1779_1), .IN6(na2966_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3265_1 ( .OUT(na3265_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2959_2), .IN6(na1781_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y74     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3266_1 ( .OUT(na3266_1), .IN1(1'b1), .IN2(~na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1783_1), .IN6(na2976_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y75     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3267_1 ( .OUT(na3267_1), .IN1(1'b1), .IN2(na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2957_2), .IN6(na1784_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a3268 ( .Y(na3268_1), .I(clk) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a3269 ( .Y(na3269_1), .I(data_in) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3270 ( .O(data_out), .A(na4154_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3271 ( .O(led[0]), .A(na4155_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3272 ( .O(led[1]), .A(na4156_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3273 ( .O(led[2]), .A(na4157_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3274 ( .O(led[3]), .A(na4158_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3275 ( .O(led[4]), .A(na4159_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3276 ( .O(led[5]), .A(na4160_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a3277 ( .Y(na3277_1), .I(reset_n) );
// C_AND///AND/      x100y99     80'h00_0078_00_0000_0C88_CCCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3278_1 ( .OUT(na3278_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2866_2), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3278_4 ( .OUT(na3278_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2802_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x144y75     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3280_2 ( .OUT(na3280_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3280_6 ( .COUTY1(na3280_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3280_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x143y96     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3281_1 ( .OUT(na3281_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1858_4), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y98     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3283_4 ( .OUT(na3283_2), .IN1(1'b1), .IN2(na2738_2), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y100     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3284_1 ( .OUT(na3284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4167_2), .IN7(1'b1), .IN8(na2071_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x121y82     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3285_4 ( .OUT(na3285_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na3151_1), .IN4(~na3150_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x113y100     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3286_1 ( .OUT(na3286_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2867_1), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3286_4 ( .OUT(na3286_2), .IN1(na15_2), .IN2(na2803_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y99     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3289_1 ( .OUT(na3289_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2739_1), .IN7(na23_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y94     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3290_4 ( .OUT(na3290_2), .IN1(na2072_1), .IN2(1'b1), .IN3(1'b1), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x109y80     80'h00_0078_00_0000_0C88_CA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3291_1 ( .OUT(na3291_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2804_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3291_4 ( .OUT(na3291_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2868_2), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y86     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3294_1 ( .OUT(na3294_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2740_1), .IN7(na23_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y91     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3295_1 ( .OUT(na3295_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4167_2), .IN7(1'b1), .IN8(na2073_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y104     80'h00_0078_00_0000_0C88_CCCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3296_1 ( .OUT(na3296_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2869_1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3296_4 ( .OUT(na3296_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2805_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y104     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3299_4 ( .OUT(na3299_2), .IN1(na2741_1), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y100     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3300_4 ( .OUT(na3300_2), .IN1(na2074_1), .IN2(1'b1), .IN3(1'b1), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y82     80'h00_0078_00_0000_0C88_AACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3301_1 ( .OUT(na3301_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(na2806_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3301_4 ( .OUT(na3301_2), .IN1(1'b1), .IN2(na2870_2), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y77     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3304_4 ( .OUT(na3304_2), .IN1(na2742_2), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y89     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3305_1 ( .OUT(na3305_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4167_2), .IN7(1'b1), .IN8(na2075_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x110y81     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3306_1 ( .OUT(na3306_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2871_1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3306_4 ( .OUT(na3306_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2807_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y71     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3309_4 ( .OUT(na3309_2), .IN1(na4171_2), .IN2(na2076_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x102y77     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3310_4 ( .OUT(na3310_2), .IN1(1'b1), .IN2(~na4167_2), .IN3(1'b1), .IN4(na2743_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y88     80'h00_0078_00_0000_0C88_F88F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3311_1 ( .OUT(na3311_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2808_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3311_4 ( .OUT(na3311_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2872_1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y89     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3314_1 ( .OUT(na3314_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na23_1), .IN8(na2424_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y85     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3315_4 ( .OUT(na3315_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2077_2), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y72     80'h00_0078_00_0000_0C88_CCCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3316_1 ( .OUT(na3316_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2873_1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3316_4 ( .OUT(na3316_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2809_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y71     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3319_1 ( .OUT(na3319_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2078_1), .IN6(na57_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y79     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3320_1 ( .OUT(na3320_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2745_2), .IN8(~na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x119y104     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3321_1 ( .OUT(na3321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2874_2), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3321_4 ( .OUT(na3321_2), .IN1(na15_2), .IN2(na2810_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y99     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3324_4 ( .OUT(na3324_2), .IN1(1'b1), .IN2(1'b1), .IN3(na23_1), .IN4(na2746_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y102     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3325_1 ( .OUT(na3325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4167_2), .IN7(1'b1), .IN8(na2079_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x132y96     80'h00_0078_00_0000_0C88_CA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3326_1 ( .OUT(na3326_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2811_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3326_4 ( .OUT(na3326_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2875_1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y97     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3329_4 ( .OUT(na3329_2), .IN1(na4166_2), .IN2(1'b1), .IN3(na2427_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y99     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3330_1 ( .OUT(na3330_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4167_2), .IN7(1'b1), .IN8(na2080_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x125y96     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3331_1 ( .OUT(na3331_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2876_2), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3331_4 ( .OUT(na3331_2), .IN1(na15_2), .IN2(na2812_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y97     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3334_4 ( .OUT(na3334_2), .IN1(1'b1), .IN2(na2748_2), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y95     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3335_4 ( .OUT(na3335_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2081_2), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x115y103     80'h00_0078_00_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3336_1 ( .OUT(na3336_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2877_1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3336_4 ( .OUT(na3336_2), .IN1(na15_2), .IN2(1'b1), .IN3(na2813_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x115y101     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3339_4 ( .OUT(na3339_2), .IN1(1'b1), .IN2(1'b1), .IN3(na23_1), .IN4(na2749_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y99     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3340_1 ( .OUT(na3340_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2082_1), .IN7(1'b1), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x125y89     80'h00_0078_00_0000_0C88_CA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3341_1 ( .OUT(na3341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2814_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3341_4 ( .OUT(na3341_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2878_2), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y94     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3344_4 ( .OUT(na3344_2), .IN1(na2750_2), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y90     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3345_4 ( .OUT(na3345_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2083_2), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x112y82     80'h00_0018_00_0000_0C88_7CFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3347_1 ( .OUT(na3347_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na103_1), .IN7(~na23_1), .IN8(~na2431_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y79     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3349_4 ( .OUT(na3349_2), .IN1(1'b1), .IN2(na4167_2), .IN3(1'b1), .IN4(na2084_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3350_1 ( .OUT(na3350_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2879_1), .IN6(~na2815_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x117y95     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3351_1 ( .OUT(na3351_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2880_2), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3351_4 ( .OUT(na3351_2), .IN1(na15_2), .IN2(1'b1), .IN3(na2816_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y97     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3354_1 ( .OUT(na3354_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2752_1), .IN7(na23_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y91     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3355_4 ( .OUT(na3355_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2085_2), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y74     80'h00_0078_00_0000_0C88_F8CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3356_1 ( .OUT(na3356_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2817_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3356_4 ( .OUT(na3356_2), .IN1(1'b1), .IN2(na2881_1), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y81     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3359_1 ( .OUT(na3359_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na23_1), .IN8(na2753_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y73     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3360_4 ( .OUT(na3360_2), .IN1(1'b1), .IN2(na4167_2), .IN3(1'b1), .IN4(na2086_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x139y108     80'h00_0078_00_0000_0C88_CCAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3361_1 ( .OUT(na3361_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2882_2), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3361_4 ( .OUT(na3361_2), .IN1(na15_2), .IN2(1'b1), .IN3(na2818_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y93     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3364_1 ( .OUT(na3364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na57_2), .IN7(na1949_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y99     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3365_1 ( .OUT(na3365_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2434_2), .IN7(1'b1), .IN8(~na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x132y94     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3366_1 ( .OUT(na3366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2883_1), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3366_4 ( .OUT(na3366_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2819_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y96     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3369_1 ( .OUT(na3369_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2435_2), .IN6(1'b1), .IN7(na23_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y96     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3370_1 ( .OUT(na3370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1950_1), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x120y99     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3371_1 ( .OUT(na3371_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2820_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3371_4 ( .OUT(na3371_2), .IN1(na2884_2), .IN2(1'b1), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x115y95     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3374_4 ( .OUT(na3374_2), .IN1(na2756_1), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y97     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3375_1 ( .OUT(na3375_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1951_2), .IN6(1'b1), .IN7(1'b1), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x122y97     80'h00_0078_00_0000_0C88_CCCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3376_1 ( .OUT(na3376_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2885_1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3376_4 ( .OUT(na3376_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2821_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y99     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3379_4 ( .OUT(na3379_2), .IN1(na2757_2), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y100     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3380_1 ( .OUT(na3380_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4167_2), .IN7(1'b1), .IN8(na1952_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x117y88     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3381_1 ( .OUT(na3381_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2886_2), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3381_4 ( .OUT(na3381_2), .IN1(na15_2), .IN2(na2822_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y88     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3384_4 ( .OUT(na3384_2), .IN1(na2758_1), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y89     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3385_1 ( .OUT(na3385_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1953_2), .IN6(1'b1), .IN7(1'b1), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x110y71     80'h00_0078_00_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3386_1 ( .OUT(na3386_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2887_1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3386_4 ( .OUT(na3386_2), .IN1(na15_2), .IN2(1'b1), .IN3(na2823_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x105y74     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3389_4 ( .OUT(na3389_2), .IN1(na2759_2), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y74     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3390_4 ( .OUT(na3390_2), .IN1(1'b1), .IN2(na4167_2), .IN3(1'b1), .IN4(na1954_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x122y82     80'h00_0078_00_0000_0C88_F88F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3391_1 ( .OUT(na3391_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2824_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3391_4 ( .OUT(na3391_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2888_2), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y88     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3394_1 ( .OUT(na3394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4166_2), .IN6(1'b1), .IN7(na2440_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y88     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3395_1 ( .OUT(na3395_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1955_2), .IN6(1'b1), .IN7(1'b1), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x104y84     80'h00_0018_00_0000_0C88_7AFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3397_1 ( .OUT(na3397_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na163_1), .IN6(1'b0), .IN7(~na23_1), .IN8(~na4335_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y78     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3399_4 ( .OUT(na3399_2), .IN1(1'b1), .IN2(na4167_2), .IN3(1'b1), .IN4(na1956_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y83     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3400_1 ( .OUT(na3400_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4310_2), .IN5(~na2825_1), .IN6(1'b0), .IN7(~na2889_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y100     80'h00_0078_00_0000_0C88_AACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3401_1 ( .OUT(na3401_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(na2826_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3401_4 ( .OUT(na3401_2), .IN1(1'b1), .IN2(na2890_2), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y98     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3404_1 ( .OUT(na3404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4166_2), .IN6(1'b1), .IN7(na2762_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y104     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3405_4 ( .OUT(na3405_2), .IN1(na3225_1), .IN2(1'b1), .IN3(1'b1), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x128y97     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3406_1 ( .OUT(na3406_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2891_1), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3406_4 ( .OUT(na3406_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2827_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y101     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3409_4 ( .OUT(na3409_2), .IN1(1'b1), .IN2(na2763_1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y97     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3410_1 ( .OUT(na3410_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3226_2), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x116y101     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3411_1 ( .OUT(na3411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2892_2), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3411_4 ( .OUT(na3411_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2828_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y102     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3414_4 ( .OUT(na3414_2), .IN1(na4166_2), .IN2(1'b1), .IN3(na2764_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y97     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3415_4 ( .OUT(na3415_2), .IN1(na3227_1), .IN2(1'b1), .IN3(1'b1), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x112y103     80'h00_0078_00_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3416_1 ( .OUT(na3416_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(na2829_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3416_4 ( .OUT(na3416_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2893_1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y99     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3419_4 ( .OUT(na3419_2), .IN1(na4166_2), .IN2(1'b1), .IN3(na2765_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y100     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3420_1 ( .OUT(na3420_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4167_2), .IN7(1'b1), .IN8(na3228_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x109y95     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3421_1 ( .OUT(na3421_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2894_2), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3421_4 ( .OUT(na3421_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2830_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x109y83     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3424_4 ( .OUT(na3424_2), .IN1(na4171_2), .IN2(na3229_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y103     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3425_4 ( .OUT(na3425_2), .IN1(1'b1), .IN2(na2766_2), .IN3(1'b1), .IN4(~na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y87     80'h00_0078_00_0000_0C88_CA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3426_1 ( .OUT(na3426_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2831_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3426_4 ( .OUT(na3426_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2895_1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y75     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3429_4 ( .OUT(na3429_2), .IN1(na4171_2), .IN2(na3230_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y91     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3430_1 ( .OUT(na3430_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2767_1), .IN7(1'b1), .IN8(~na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x109y94     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3431_1 ( .OUT(na3431_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2896_2), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3431_4 ( .OUT(na3431_2), .IN1(na15_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2832_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y96     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3434_4 ( .OUT(na3434_2), .IN1(1'b1), .IN2(na2768_2), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y92     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3435_1 ( .OUT(na3435_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3231_1), .IN7(1'b1), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y90     80'h00_0078_00_0000_0C88_CACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3436_1 ( .OUT(na3436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2833_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3436_4 ( .OUT(na3436_2), .IN1(1'b1), .IN2(na2897_1), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y99     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3439_1 ( .OUT(na3439_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2769_1), .IN6(1'b1), .IN7(na23_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y87     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3440_4 ( .OUT(na3440_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3232_2), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y111     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3441_1 ( .OUT(na3441_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na241_1), .IN7(na240_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x121y113     80'h00_0060_00_0000_0C06_FFC3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3442_4 ( .OUT(na3442_2), .IN1(1'b0), .IN2(~na1797_1), .IN3(1'b0), .IN4(na1801_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y111     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3446_1 ( .OUT(na3446_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3010_2), .IN6(1'b0), .IN7(1'b0), .IN8(na227_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x125y116     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3447_1 ( .OUT(na3447_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na223_1), .IN6(1'b0), .IN7(1'b0), .IN8(na227_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x128y113     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3449_4 ( .OUT(na3449_2), .IN1(na226_1), .IN2(1'b0), .IN3(1'b0), .IN4(na230_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y115     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3451_1 ( .OUT(na3451_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1797_1), .IN7(na1799_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y111     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3452_4 ( .OUT(na3452_2), .IN1(1'b0), .IN2(1'b0), .IN3(na246_1), .IN4(~na248_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y113     80'h00_0018_00_0000_0C66_C300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3453_1 ( .OUT(na3453_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na232_1), .IN7(1'b0), .IN8(na1801_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y115     80'h00_0060_00_0000_0C06_FF53
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3454_4 ( .OUT(na3454_2), .IN1(1'b0), .IN2(~na232_1), .IN3(~na1799_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y109     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3455_1 ( .OUT(na3455_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na226_1), .IN6(na244_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x127y112     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3456_4 ( .OUT(na3456_2), .IN1(na220_2), .IN2(1'b0), .IN3(na222_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y113     80'h00_0060_00_0000_0C06_FFA3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3457_4 ( .OUT(na3457_2), .IN1(1'b0), .IN2(~na253_2), .IN3(na242_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y107     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3462_1 ( .OUT(na3462_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3010_2), .IN6(na244_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y107     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3463_4 ( .OUT(na3463_2), .IN1(1'b0), .IN2(1'b0), .IN3(na240_2), .IN4(~na248_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y83     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3465_1 ( .OUT(na3465_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na57_2), .IN7(na2087_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y91     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3466_1 ( .OUT(na3466_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2906_2), .IN7(1'b1), .IN8(~na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x128y112     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3470_1 ( .OUT(na3470_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na247_2), .IN7(na240_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y108     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3472_4 ( .OUT(na3472_2), .IN1(1'b0), .IN2(na241_1), .IN3(na246_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y88     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3474_1 ( .OUT(na3474_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4171_2), .IN6(na2088_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y94     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3475_4 ( .OUT(na3475_2), .IN1(na2907_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y81     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3479_1 ( .OUT(na3479_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na57_2), .IN7(1'b1), .IN8(na2089_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y81     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3480_4 ( .OUT(na3480_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2908_2), .IN4(~na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x131y111     80'h00_0060_00_0000_0C06_FF5C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3483_4 ( .OUT(na3483_2), .IN1(1'b0), .IN2(na253_2), .IN3(~na222_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x128y111     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3484_1 ( .OUT(na3484_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na220_2), .IN6(1'b0), .IN7(na242_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x117y90     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3486_1 ( .OUT(na3486_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3489_1), .IN6(~na16_2), .IN7(1'b0), .IN8(~na290_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y91     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3489_1 ( .OUT(na3489_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2409_1), .IN8(~na2322_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x113y92     80'h00_0060_00_0000_0C08_FF7C
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3490_4 ( .OUT(na3490_2), .IN1(1'b0), .IN2(na292_1), .IN3(~na23_1), .IN4(~na2909_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y96     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3492_4 ( .OUT(na3492_2), .IN1(1'b1), .IN2(na4167_2), .IN3(1'b1), .IN4(na2090_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y75     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3494_1 ( .OUT(na3494_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na57_2), .IN7(1'b1), .IN8(na2091_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y79     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3495_4 ( .OUT(na3495_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2910_2), .IN4(~na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x113y79     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3499_1 ( .OUT(na3499_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3502_1), .IN6(~na16_2), .IN7(1'b0), .IN8(~na305_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x117y83     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3502_1 ( .OUT(na3502_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2411_1), .IN6(1'b0), .IN7(~na2324_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y70     80'h00_0018_00_0000_0C88_C7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3503_1 ( .OUT(na3503_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2092_1), .IN6(~na57_2), .IN7(1'b0), .IN8(na307_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x103y81     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3505_4 ( .OUT(na3505_2), .IN1(na2911_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x110y82     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3507_4 ( .OUT(na3507_2), .IN1(1'b1), .IN2(na2912_2), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y87     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3508_1 ( .OUT(na3508_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2093_2), .IN8(na24_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y84     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3512_1 ( .OUT(na3512_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2913_1), .IN7(na23_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y74     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3513_4 ( .OUT(na3513_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2094_1), .IN4(na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x140y81     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3516_1 ( .OUT(na3516_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na323_2), .IN6(na3002_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x132y86     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3518_4 ( .OUT(na3518_2), .IN1(~na15_2), .IN2(~na2351_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x139y83     80'h00_0078_00_0000_0C88_8F8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3519_1 ( .OUT(na3519_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na322_1), .IN8(na2311_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3519_4 ( .OUT(na3519_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2978_2), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y84     80'h00_0018_00_0000_0888_1F34
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3523_1 ( .OUT(na3523_1), .IN1(~na334_1), .IN2(na332_1), .IN3(1'b1), .IN4(~na3528_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na335_1),
                      .IN8(~na3528_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x140y86     80'h00_0078_00_0000_0C88_CA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3528_1 ( .OUT(na3528_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na323_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3003_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3528_4 ( .OUT(na3528_2), .IN1(1'b1), .IN2(1'b1), .IN3(na322_1), .IN4(na2312_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y95     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3529_1 ( .OUT(na3529_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2979_1), .IN8(~na2352_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y79     80'h00_0018_00_0000_0888_4513
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3531_1 ( .OUT(na3531_1), .IN1(1'b1), .IN2(~na344_1), .IN3(~na3534_1), .IN4(~na3532_1), .IN5(~na343_1), .IN6(1'b1), .IN7(~na3534_2),
                      .IN8(na3533_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y86     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3532_1 ( .OUT(na3532_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2353_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x138y78     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3533_4 ( .OUT(na3533_2), .IN1(~na2980_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x142y79     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3534_1 ( .OUT(na3534_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2313_1), .IN8(na4192_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3534_4 ( .OUT(na3534_2), .IN1(na323_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3004_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y82     80'h00_0018_00_0000_0888_5145
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3540_1 ( .OUT(na3540_1), .IN1(~na353_1), .IN2(1'b1), .IN3(~na3543_1), .IN4(na3542_1), .IN5(~na3541_1), .IN6(~na352_1), .IN7(~na3543_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y79     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3541_1 ( .OUT(na3541_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3005_1), .IN6(1'b1), .IN7(na4194_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x126y86     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3542_1 ( .OUT(na3542_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na15_2), .IN6(1'b0), .IN7(~na2354_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x136y81     80'h00_0078_00_0000_0C88_8F8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3543_1 ( .OUT(na3543_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na322_1), .IN8(na2314_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3543_4 ( .OUT(na3543_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2981_1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x140y68     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3548_4 ( .OUT(na3548_2), .IN1(1'b1), .IN2(na2315_1), .IN3(na322_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x133y74     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3550_4 ( .OUT(na3550_2), .IN1(~na15_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na2355_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x138y73     80'h00_0078_00_0000_0C88_CACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3551_1 ( .OUT(na3551_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na323_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3006_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3551_4 ( .OUT(na3551_2), .IN1(1'b1), .IN2(na2982_2), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y69     80'h00_0018_00_0000_0888_5541
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3555_1 ( .OUT(na3555_1), .IN1(~na3556_1), .IN2(~na371_1), .IN3(~na3558_1), .IN4(na3557_2), .IN5(~na370_1), .IN6(1'b1), .IN7(~na3558_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x127y75     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3556_1 ( .OUT(na3556_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2356_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x134y72     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3557_4 ( .OUT(na3557_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na2983_1), .IN4(~na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x136y69     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3558_1 ( .OUT(na3558_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2316_2), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3558_4 ( .OUT(na3558_2), .IN1(na323_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3007_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x136y75     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3563_1 ( .OUT(na3563_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3008_2), .IN6(na4195_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x130y82     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3565_1 ( .OUT(na3565_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na15_2), .IN6(~na2357_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x137y77     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3566_1 ( .OUT(na3566_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2317_1), .IN6(1'b1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3566_4 ( .OUT(na3566_2), .IN1(na2984_2), .IN2(1'b1), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x134y69     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3570_1 ( .OUT(na3570_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2318_2), .IN8(na4192_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3570_4 ( .OUT(na3570_2), .IN1(na323_2), .IN2(na3009_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y79     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3572_1 ( .OUT(na3572_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2985_1), .IN6(~na2358_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x109y93     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3576_1 ( .OUT(na3576_1), .IN1(na21_2), .IN2(~na2055_2), .IN3(~na1991_1), .IN4(na19_1), .IN5(~na2023_2), .IN6(~na16_2), .IN7(na26_2),
                      .IN8(~na1959_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y84     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3577_4 ( .OUT(na3577_2), .IN1(na3042_2), .IN2(na4195_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x134y91     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3579_1 ( .OUT(na3579_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na15_2), .IN6(1'b0), .IN7(~na2383_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x139y86     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3580_1 ( .OUT(na3580_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2343_1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3580_4 ( .OUT(na3580_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2986_2), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x136y87     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3585_1 ( .OUT(na3585_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2987_2), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3585_4 ( .OUT(na3585_2), .IN1(na15_2), .IN2(1'b1), .IN3(na2384_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x140y70     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3590_4 ( .OUT(na3590_2), .IN1(1'b1), .IN2(na4193_2), .IN3(na2345_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x136y77     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3592_1 ( .OUT(na3592_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2988_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x137y76     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3593_1 ( .OUT(na3593_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na323_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3044_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3593_4 ( .OUT(na3593_2), .IN1(na15_2), .IN2(na2385_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x141y82     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3597_4 ( .OUT(na3597_2), .IN1(na2989_1), .IN2(1'b1), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x135y83     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3598_1 ( .OUT(na3598_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na15_2), .IN6(~na2386_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x140y80     80'h00_0078_00_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3599_1 ( .OUT(na3599_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3045_1), .IN6(1'b1), .IN7(na4194_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3599_4 ( .OUT(na3599_2), .IN1(1'b1), .IN2(1'b1), .IN3(na322_1), .IN4(na2346_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y69     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3604_4 ( .OUT(na3604_2), .IN1(na323_2), .IN2(na3046_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x131y72     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3606_1 ( .OUT(na3606_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na15_2), .IN6(~na2387_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x133y69     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3607_1 ( .OUT(na3607_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2347_1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3607_4 ( .OUT(na3607_2), .IN1(1'b1), .IN2(1'b1), .IN3(na4169_2), .IN4(na2990_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y77     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3611_1 ( .OUT(na3611_1), .IN1(na21_2), .IN2(~na2060_1), .IN3(~na1996_1), .IN4(na19_1), .IN5(~na2028_1), .IN6(~na16_2), .IN7(na26_2),
                      .IN8(~na1964_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x136y68     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3612_1 ( .OUT(na3612_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na323_2), .IN6(1'b1), .IN7(na3047_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x130y71     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3614_4 ( .OUT(na3614_2), .IN1(~na15_2), .IN2(~na2388_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x135y66     80'h00_0078_00_0000_0C88_8F8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3615_1 ( .OUT(na3615_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2348_2), .IN8(na4192_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3615_4 ( .OUT(na3615_2), .IN1(1'b1), .IN2(1'b1), .IN3(na4169_2), .IN4(na2991_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x135y74     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3620_1 ( .OUT(na3620_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2992_2), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x134y73     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3621_4 ( .OUT(na3621_2), .IN1(~na15_2), .IN2(1'b0), .IN3(~na2389_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x138y72     80'h00_0078_00_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3622_1 ( .OUT(na3622_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3048_2), .IN6(1'b1), .IN7(na4194_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3622_4 ( .OUT(na3622_2), .IN1(1'b1), .IN2(na2349_1), .IN3(na322_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x135y67     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3627_1 ( .OUT(na3627_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2350_2), .IN6(1'b1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3627_4 ( .OUT(na3627_2), .IN1(na323_2), .IN2(na3049_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y75     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3629_1 ( .OUT(na3629_1), .IN1(1'b1), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2993_1), .IN8(~na2390_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x131y86     80'h00_0018_00_0000_0888_3512
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3633_1 ( .OUT(na3633_1), .IN1(na3635_2), .IN2(~na468_1), .IN3(~na3634_1), .IN4(~na3636_1), .IN5(~na467_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na3636_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y91     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3634_1 ( .OUT(na3634_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2914_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x133y87     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3635_4 ( .OUT(na3635_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na3050_2), .IN4(~na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x136y86     80'h00_0078_00_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3636_1 ( .OUT(na3636_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na323_2), .IN6(1'b1), .IN7(na3058_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3636_4 ( .OUT(na3636_2), .IN1(1'b1), .IN2(na2375_1), .IN3(na322_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x117y93     80'h00_0018_00_0000_0888_B7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3641_1 ( .OUT(na3641_1), .IN1(na21_2), .IN2(~na2048_1), .IN3(~na1984_1), .IN4(na19_1), .IN5(~na2016_1), .IN6(~na16_2), .IN7(na26_2),
                      .IN8(~na3187_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y87     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3642_1 ( .OUT(na3642_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3051_1), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x139y96     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3643_4 ( .OUT(na3643_2), .IN1(~na15_2), .IN2(1'b0), .IN3(~na2915_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x138y88     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3644_1 ( .OUT(na3644_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2376_2), .IN8(na4192_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3644_4 ( .OUT(na3644_2), .IN1(na323_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3059_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y80     80'h00_0018_00_0000_0888_3512
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3650_1 ( .OUT(na3650_1), .IN1(na3652_2), .IN2(~na485_1), .IN3(~na3651_1), .IN4(~na3653_1), .IN5(~na484_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na3653_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y85     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3651_1 ( .OUT(na3651_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(1'b1), .IN7(na2916_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x135y83     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3652_4 ( .OUT(na3652_2), .IN1(~na3052_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x138y80     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3653_1 ( .OUT(na3653_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2377_1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3653_4 ( .OUT(na3653_2), .IN1(na323_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3060_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x122y86     80'h00_0018_00_0000_0888_A313
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3659_1 ( .OUT(na3659_1), .IN1(1'b1), .IN2(~na494_1), .IN3(~na4398_2), .IN4(~na493_1), .IN5(1'b1), .IN6(~na3663_2), .IN7(na491_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x123y84     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3663_1 ( .OUT(na3663_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_2), .IN6(na2917_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3663_4 ( .OUT(na3663_2), .IN1(na3053_1), .IN2(1'b1), .IN3(1'b1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y77     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3665_1 ( .OUT(na3665_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3062_2), .IN6(na4195_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x135y78     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3667_4 ( .OUT(na3667_2), .IN1(~na15_2), .IN2(1'b0), .IN3(~na2918_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x139y73     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3668_1 ( .OUT(na3668_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2379_1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3668_4 ( .OUT(na3668_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3054_1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y70     80'h00_0018_00_0000_0888_5312
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3672_1 ( .OUT(na3672_1), .IN1(na3674_1), .IN2(~na3673_1), .IN3(~na3675_1), .IN4(~na509_1), .IN5(1'b1), .IN6(~na508_1), .IN7(~na3675_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x137y74     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3673_1 ( .OUT(na3673_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3063_1), .IN6(na4195_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x127y77     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3674_1 ( .OUT(na3674_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na15_2), .IN6(1'b0), .IN7(~na2919_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x132y73     80'h00_0078_00_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3675_1 ( .OUT(na3675_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2380_2), .IN6(1'b1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3675_4 ( .OUT(na3675_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3055_1), .IN4(na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y80     80'h00_0018_00_0000_0888_1F12
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3680_1 ( .OUT(na3680_1), .IN1(na3682_1), .IN2(~na521_1), .IN3(~na3683_1), .IN4(~na3681_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na3683_2),
                      .IN8(~na520_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y86     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3681_4 ( .OUT(na3681_2), .IN1(na15_2), .IN2(na2920_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x127y81     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3682_1 ( .OUT(na3682_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na3056_2), .IN8(~na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x130y81     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3683_1 ( .OUT(na3683_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2381_1), .IN6(1'b1), .IN7(na322_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3683_4 ( .OUT(na3683_2), .IN1(na323_2), .IN2(na3064_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x125y81     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3689_1 ( .OUT(na3689_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3057_1), .IN6(1'b1), .IN7(1'b1), .IN8(na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3689_4 ( .OUT(na3689_2), .IN1(na15_2), .IN2(1'b1), .IN3(na2921_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y72     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3694_4 ( .OUT(na3694_2), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(~na3150_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y74     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3695_1 ( .OUT(na3695_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na539_2), .IN7(~na1947_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x139y66     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3696_1 ( .OUT(na3696_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na533_1), .IN6(na1957_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y111     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3699_4 ( .OUT(na3699_2), .IN1(1'b0), .IN2(na830_1), .IN3(na815_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y115     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3700_1 ( .OUT(na3700_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na824_1), .IN8(na1836_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x144y112     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3704_4 ( .OUT(na3704_2), .IN1(na3025_2), .IN2(1'b0), .IN3(na3019_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x149y116     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3705_1 ( .OUT(na3705_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na813_1), .IN7(na812_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y113     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3707_4 ( .OUT(na3707_2), .IN1(na814_1), .IN2(1'b1), .IN3(~na812_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y116     80'h00_0018_00_0000_0C66_5C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3709_1 ( .OUT(na3709_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na813_1), .IN7(~na3018_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y113     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3711_1 ( .OUT(na3711_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na819_1), .IN7(1'b0), .IN8(na1836_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x144y109     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3712_4 ( .OUT(na3712_2), .IN1(na814_1), .IN2(na818_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y114     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3713_1 ( .OUT(na3713_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1834_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1836_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y116     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3714_4 ( .OUT(na3714_2), .IN1(na1834_1), .IN2(1'b0), .IN3(~na824_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y107     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3716_1 ( .OUT(na3716_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na836_2), .IN8(na837_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x142y107     80'h00_0078_00_0000_0C88_F853
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3717_1 ( .OUT(na3717_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na814_1), .IN6(na830_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3717_4 ( .OUT(na3717_2), .IN1(1'b1), .IN2(~na818_1), .IN3(~na832_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y111     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3720_1 ( .OUT(na3720_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na843_1), .IN6(1'b0), .IN7(na842_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y109     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3721_1 ( .OUT(na3721_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na847_1), .IN6(1'b0), .IN7(1'b0), .IN8(na845_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x142y112     80'h00_0060_00_0000_0C06_FF5C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3722_4 ( .OUT(na3722_2), .IN1(1'b0), .IN2(na830_1), .IN3(~na3018_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x142y112     80'h00_0018_00_0000_0C66_5A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3723_1 ( .OUT(na3723_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na847_1), .IN6(1'b0), .IN7(~na842_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x130y91     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3724_1 ( .OUT(na3724_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3244_1), .IN6(1'b0), .IN7(na3106_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x147y116     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3726_4 ( .OUT(na3726_2), .IN1(na843_1), .IN2(1'b0), .IN3(1'b0), .IN4(na845_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y109     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3728_4 ( .OUT(na3728_2), .IN1(1'b0), .IN2(na846_1), .IN3(na842_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y98     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3729_4 ( .OUT(na3729_2), .IN1(1'b0), .IN2(na3107_1), .IN3(1'b0), .IN4(na3245_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y85     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3730_1 ( .OUT(na3730_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3108_2), .IN6(na3246_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y108     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3731_4 ( .OUT(na3731_2), .IN1(1'b0), .IN2(na818_1), .IN3(na836_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y105     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3732_1 ( .OUT(na3732_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na814_1), .IN6(1'b0), .IN7(1'b0), .IN8(na837_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y90     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3733_1 ( .OUT(na3733_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3247_1), .IN8(na3109_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x132y75     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3734_4 ( .OUT(na3734_2), .IN1(na3248_1), .IN2(1'b0), .IN3(na3110_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y76     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3735_1 ( .OUT(na3735_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3249_1), .IN8(na3111_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x133y86     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3736_4 ( .OUT(na3736_2), .IN1(na3112_2), .IN2(na3250_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x128y76     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3737_1 ( .OUT(na3737_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3113_2), .IN8(na3251_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y106     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3738_4 ( .OUT(na3738_2), .IN1(na903_1), .IN2(1'b0), .IN3(~na3026_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x149y105     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3739_1 ( .OUT(na3739_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1843_2), .IN7(1'b0), .IN8(na1841_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x149y109     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3741_4 ( .OUT(na3741_2), .IN1(1'b1), .IN2(na894_2), .IN3(~na897_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y99     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3742_1 ( .OUT(na3742_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3027_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na3033_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x147y104     80'h00_0060_00_0000_0C06_FFC9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3744_4 ( .OUT(na3744_2), .IN1(na3027_1), .IN2(~na4370_2), .IN3(1'b0), .IN4(na891_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x149y102     80'h00_0060_00_0000_0C06_FF35
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3748_4 ( .OUT(na3748_2), .IN1(~na3027_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na3033_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x150y102     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3749_1 ( .OUT(na3749_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1839_1), .IN6(na1843_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x148y100     80'h00_0060_00_0000_0C06_FFA5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3750_4 ( .OUT(na3750_2), .IN1(~na908_1), .IN2(1'b0), .IN3(na909_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y102     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3751_1 ( .OUT(na3751_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1839_1), .IN6(1'b0), .IN7(na888_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x147y106     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3752_4 ( .OUT(na3752_2), .IN1(1'b0), .IN2(1'b0), .IN3(na888_1), .IN4(na1841_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y99     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3756_1 ( .OUT(na3756_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na908_1), .IN6(1'b0), .IN7(1'b0), .IN8(na907_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y97     80'h00_0060_00_0000_0C06_FF5C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3757_4 ( .OUT(na3757_2), .IN1(1'b0), .IN2(na918_2), .IN3(~na909_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y104     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3758_1 ( .OUT(na3758_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na903_1), .IN6(1'b0), .IN7(1'b0), .IN8(na893_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x144y105     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3759_4 ( .OUT(na3759_2), .IN1(~na892_2), .IN2(1'b0), .IN3(1'b0), .IN4(na907_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y99     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3760_1 ( .OUT(na3760_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na887_1), .IN7(1'b0), .IN8(na907_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x144y103     80'h00_0060_00_0000_0C06_FFC3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3761_4 ( .OUT(na3761_2), .IN1(1'b0), .IN2(~na924_1), .IN3(1'b0), .IN4(na916_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x136y93     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3762_4 ( .OUT(na3762_2), .IN1(na3114_2), .IN2(1'b0), .IN3(1'b0), .IN4(na3252_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y98     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3764_1 ( .OUT(na3764_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na908_1), .IN6(1'b0), .IN7(1'b0), .IN8(na904_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x148y102     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3766_4 ( .OUT(na3766_2), .IN1(1'b0), .IN2(na918_2), .IN3(na915_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x140y91     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3767_4 ( .OUT(na3767_2), .IN1(1'b0), .IN2(na3253_1), .IN3(na3115_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y81     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3768_1 ( .OUT(na3768_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3254_1), .IN6(1'b0), .IN7(na3116_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y103     80'h00_0060_00_0000_0C06_FF5C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3769_4 ( .OUT(na3769_2), .IN1(1'b0), .IN2(na924_1), .IN3(~na897_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y103     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3770_4 ( .OUT(na3770_2), .IN1(~na892_2), .IN2(1'b0), .IN3(1'b0), .IN4(na916_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x132y90     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3771_1 ( .OUT(na3771_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3255_1), .IN7(1'b0), .IN8(na3117_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x130y75     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3772_1 ( .OUT(na3772_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3256_1), .IN7(na3118_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y70     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3773_4 ( .OUT(na3773_2), .IN1(na3119_1), .IN2(na3257_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y69     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3774_4 ( .OUT(na3774_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3120_2), .IN4(na3258_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y72     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3775_1 ( .OUT(na3775_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3259_1), .IN8(na3121_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x136y113     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3778_4 ( .OUT(na3778_2), .IN1(1'b0), .IN2(na970_1), .IN3(1'b0), .IN4(na1848_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y114     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3781_1 ( .OUT(na3781_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3035_1), .IN7(1'b0), .IN8(na3041_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y117     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3782_4 ( .OUT(na3782_2), .IN1(1'b0), .IN2(na964_1), .IN3(na965_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y115     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3784_1 ( .OUT(na3784_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na963_2), .IN6(1'b1), .IN7(~na965_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x139y116     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3785_4 ( .OUT(na3785_2), .IN1(na3034_2), .IN2(1'b0), .IN3(1'b0), .IN4(na969_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x133y115     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3788_4 ( .OUT(na3788_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1846_2), .IN4(na1848_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y115     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3790_1 ( .OUT(na3790_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na975_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1848_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x137y116     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3792_4 ( .OUT(na3792_2), .IN1(na975_1), .IN2(1'b0), .IN3(na1846_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y113     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3794_1 ( .OUT(na3794_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na988_1), .IN6(1'b0), .IN7(na989_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y115     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3795_1 ( .OUT(na3795_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na988_1), .IN6(na984_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x132y114     80'h00_0060_00_0000_0C06_FF5C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3796_4 ( .OUT(na3796_2), .IN1(1'b0), .IN2(na995_2), .IN3(~na989_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y116     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3798_1 ( .OUT(na3798_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na963_2), .IN6(na984_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x132y115     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3799_4 ( .OUT(na3799_2), .IN1(1'b0), .IN2(na984_1), .IN3(1'b0), .IN4(na983_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x132y113     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3800_1 ( .OUT(na3800_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1001_2), .IN6(1'b0), .IN7(1'b0), .IN8(na993_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x135y94     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3801_4 ( .OUT(na3801_2), .IN1(1'b0), .IN2(na3122_2), .IN3(1'b0), .IN4(na3260_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x130y116     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3803_1 ( .OUT(na3803_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na995_2), .IN7(na992_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x130y115     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3805_4 ( .OUT(na3805_2), .IN1(na988_1), .IN2(1'b0), .IN3(1'b0), .IN4(na986_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y95     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3806_1 ( .OUT(na3806_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3123_1), .IN7(na3261_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x135y90     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3807_4 ( .OUT(na3807_2), .IN1(1'b0), .IN2(na3262_1), .IN3(na3124_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x133y112     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3808_1 ( .OUT(na3808_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1001_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na969_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x135y114     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3809_4 ( .OUT(na3809_2), .IN1(~na963_2), .IN2(1'b0), .IN3(1'b0), .IN4(na993_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y91     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3810_1 ( .OUT(na3810_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3263_1), .IN7(1'b0), .IN8(na3125_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x135y88     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3811_4 ( .OUT(na3811_2), .IN1(na3126_2), .IN2(1'b0), .IN3(1'b0), .IN4(na3264_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y77     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3812_1 ( .OUT(na3812_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3265_1), .IN7(1'b0), .IN8(na3127_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x128y89     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3813_4 ( .OUT(na3813_2), .IN1(1'b0), .IN2(na3266_1), .IN3(na3128_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y83     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3814_1 ( .OUT(na3814_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3267_1), .IN6(na3129_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x124y84     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3863_4 ( .OUT(na3863_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3236_1), .IN4(na3098_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y91     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3864_1 ( .OUT(na3864_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3099_1), .IN7(1'b0), .IN8(na3237_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y75     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3865_4 ( .OUT(na3865_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3100_2), .IN4(na3238_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y91     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3866_1 ( .OUT(na3866_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3101_1), .IN7(1'b0), .IN8(na3239_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x119y73     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3867_4 ( .OUT(na3867_2), .IN1(1'b0), .IN2(na3240_1), .IN3(1'b0), .IN4(na3102_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y80     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3868_1 ( .OUT(na3868_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3241_1), .IN7(na3103_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y81     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3869_1 ( .OUT(na3869_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3242_1), .IN7(1'b0), .IN8(na3104_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y76     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3870_4 ( .OUT(na3870_2), .IN1(na3243_1), .IN2(1'b0), .IN3(1'b0), .IN4(na3105_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y90     80'h00_0018_00_0000_0888_AC12
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3944_1 ( .OUT(na3944_1), .IN1(na1217_1), .IN2(~na1214_1), .IN3(~na3948_1), .IN4(~na3946_2), .IN5(1'b1), .IN6(na3947_1), .IN7(na3945_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x142y85     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3945_1 ( .OUT(na3945_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1206_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na2406_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y88     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3946_4 ( .OUT(na3946_2), .IN1(na3074_2), .IN2(1'b1), .IN3(na1208_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x141y86     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3947_1 ( .OUT(na3947_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1211_2), .IN6(1'b0), .IN7(~na3134_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y87     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3948_1 ( .OUT(na3948_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2994_2), .IN6(1'b1), .IN7(na1212_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y95     80'h00_0018_00_0000_0888_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3950_1 ( .OUT(na3950_1), .IN1(~na1945_2), .IN2(~na4301_2), .IN3(~na1943_1), .IN4(~na1946_1), .IN5(~na1945_1), .IN6(~na1941_2),
                      .IN7(~na4300_2), .IN8(~na1946_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x140y82     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3951_1 ( .OUT(na3951_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1219_2), .IN6(1'b0), .IN7(~na2898_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x143y85     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3952_1 ( .OUT(na3952_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3002_2), .IN7(na1220_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x147y86     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3953_4 ( .OUT(na3953_2), .IN1(~na3042_2), .IN2(1'b0), .IN3(~na1222_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x143y88     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3954_4 ( .OUT(na3954_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3058_2), .IN4(na4264_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x145y87     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3955_1 ( .OUT(na3955_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1226_2), .IN7(~na2986_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y87     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3956_4 ( .OUT(na3956_2), .IN1(1'b1), .IN2(na1227_1), .IN3(na3050_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x142y91     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3957_1 ( .OUT(na3957_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2938_2), .IN6(~na1229_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y90     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3958_1 ( .OUT(na3958_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3090_2), .IN8(na1230_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x144y91     80'h00_0078_00_0000_0CEE_3553
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3959_1 ( .OUT(na3959_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1232_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na3066_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3959_4 ( .OUT(na3959_2), .IN1(1'b0), .IN2(~na1920_1), .IN3(~na1235_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y90     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3960_4 ( .OUT(na3960_2), .IN1(1'b1), .IN2(na3082_2), .IN3(1'b1), .IN4(na1233_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y88     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3962_1 ( .OUT(na3962_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2978_2), .IN8(na1236_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y91     80'h00_0018_00_0000_0888_8841
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3963_1 ( .OUT(na3963_1), .IN1(~na1239_1), .IN2(~na3966_2), .IN3(~na3964_2), .IN4(na1242_2), .IN5(na1243_1), .IN6(na3965_1),
                      .IN7(na1244_1), .IN8(na1245_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y89     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3964_4 ( .OUT(na3964_2), .IN1(na3051_1), .IN2(na1227_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x141y92     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3965_1 ( .OUT(na3965_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1921_2), .IN6(1'b0), .IN7(~na1235_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x141y88     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3966_4 ( .OUT(na3966_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2979_1), .IN4(na1236_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x142y89     80'h00_0078_00_0000_0CEE_5335
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3975_1 ( .OUT(na3975_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3075_1), .IN7(~na1208_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3975_4 ( .OUT(na3975_2), .IN1(~na1211_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na3135_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y86     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3976_4 ( .OUT(na3976_2), .IN1(na2987_2), .IN2(na1226_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y87     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3978_4 ( .OUT(na3978_2), .IN1(na4263_2), .IN2(1'b1), .IN3(na3043_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y81     80'h00_0018_00_0000_0888_4242
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3979_1 ( .OUT(na3979_1), .IN1(na1255_1), .IN2(~na1251_2), .IN3(~na3984_1), .IN4(na1254_1), .IN5(na3981_2), .IN6(~na3980_1),
                      .IN7(~na3984_2), .IN8(na3983_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y80     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3980_1 ( .OUT(na3980_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1222_2), .IN8(na3044_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x143y81     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3981_4 ( .OUT(na3981_2), .IN1(~na1232_1), .IN2(1'b0), .IN3(~na3068_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x146y84     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3983_1 ( .OUT(na3983_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3076_2), .IN6(1'b0), .IN7(~na1208_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x144y83     80'h00_0078_00_0000_0C88_8FCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3984_1 ( .OUT(na3984_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3084_2), .IN8(na1233_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3984_4 ( .OUT(na3984_2), .IN1(1'b1), .IN2(na1229_2), .IN3(1'b1), .IN4(na2940_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x142y81     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3990_1 ( .OUT(na3990_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1211_2), .IN6(~na3136_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3990_4 ( .OUT(na3990_2), .IN1(~na1206_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na2408_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y82     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3991_1 ( .OUT(na3991_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1220_1), .IN8(na3004_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y85     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3993_1 ( .OUT(na3993_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1224_2), .IN8(na3060_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y87     80'h00_0018_00_0000_0888_8814
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3994_1 ( .OUT(na3994_1), .IN1(~na3997_2), .IN2(na1265_2), .IN3(~na3995_2), .IN4(~na1262_2), .IN5(na1266_1), .IN6(na1268_2),
                      .IN7(na3996_1), .IN8(na1267_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x140y85     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3995_4 ( .OUT(na3995_2), .IN1(na1206_2), .IN2(1'b1), .IN3(na2409_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x142y87     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3996_1 ( .OUT(na3996_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2997_1), .IN6(1'b0), .IN7(~na1212_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x141y87     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3997_4 ( .OUT(na3997_2), .IN1(na2941_1), .IN2(na1229_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x143y89     80'h00_0078_00_0000_0CEE_7007
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4006_1 ( .OUT(na4006_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na3085_1), .IN8(~na1233_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4006_4 ( .OUT(na4006_2), .IN1(~na1232_1), .IN2(~na3069_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y86     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4007_4 ( .OUT(na4007_2), .IN1(na3045_1), .IN2(1'b1), .IN3(na1222_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y90     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4009_1 ( .OUT(na4009_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3061_1), .IN6(1'b1), .IN7(na1224_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x141y78     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4010_1 ( .OUT(na4010_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1211_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na3138_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y78     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4011_1 ( .OUT(na4011_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1227_1), .IN7(na3054_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x143y77     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4012_1 ( .OUT(na4012_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3086_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na1233_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y81     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4013_1 ( .OUT(na4013_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3094_2), .IN7(1'b1), .IN8(na1230_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x142y75     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4014_1 ( .OUT(na4014_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2410_2), .IN6(1'b0), .IN7(~na4259_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y78     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4015_4 ( .OUT(na4015_2), .IN1(na3070_2), .IN2(na4265_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x143y79     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4018_1 ( .OUT(na4018_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3078_2), .IN6(1'b0), .IN7(~na1208_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x140y78     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4019_4 ( .OUT(na4019_2), .IN1(1'b1), .IN2(na1924_1), .IN3(na1235_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x147y78     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4020_1 ( .OUT(na4020_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na2982_2), .IN7(1'b0), .IN8(~na1236_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y73     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4021_4 ( .OUT(na4021_2), .IN1(1'b1), .IN2(na1226_2), .IN3(1'b1), .IN4(na2990_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x144y78     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4022_1 ( .OUT(na4022_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2998_2), .IN6(1'b0), .IN7(~na1212_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y79     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4023_4 ( .OUT(na4023_2), .IN1(na3062_2), .IN2(1'b1), .IN3(na1224_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x140y77     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4024_1 ( .OUT(na4024_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1219_2), .IN6(~na2902_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y82     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4025_4 ( .OUT(na4025_2), .IN1(1'b1), .IN2(na1229_2), .IN3(na2942_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x141y72     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4026_1 ( .OUT(na4026_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1226_2), .IN7(1'b0), .IN8(~na2991_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x143y78     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4027_4 ( .OUT(na4027_2), .IN1(1'b1), .IN2(na3095_1), .IN3(1'b1), .IN4(na1230_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x140y71     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4028_1 ( .OUT(na4028_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1211_2), .IN6(~na3139_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x141y73     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4029_4 ( .OUT(na4029_2), .IN1(na3087_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1233_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x142y78     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4030_1 ( .OUT(na4030_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na2999_1), .IN7(~na1212_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x142y76     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4031_4 ( .OUT(na4031_2), .IN1(na1219_2), .IN2(1'b1), .IN3(na2903_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x143y75     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4034_1 ( .OUT(na4034_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1220_1), .IN8(~na3007_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y73     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4035_4 ( .OUT(na4035_2), .IN1(1'b1), .IN2(na1227_1), .IN3(na3055_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x141y76     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4036_4 ( .OUT(na4036_2), .IN1(~na2411_1), .IN2(1'b0), .IN3(~na4259_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x142y73     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4037_1 ( .OUT(na4037_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1232_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3071_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x142y70     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4038_4 ( .OUT(na4038_2), .IN1(~na4263_2), .IN2(1'b0), .IN3(~na3047_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x143y76     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4039_1 ( .OUT(na4039_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3063_1), .IN6(1'b1), .IN7(na1224_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x142y75     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4040_4 ( .OUT(na4040_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1208_1), .IN4(~na3079_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x140y78     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4041_1 ( .OUT(na4041_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1235_1), .IN8(na1925_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y79     80'h00_0018_00_0000_0888_8814
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4042_1 ( .OUT(na4042_1), .IN1(~na1295_1), .IN2(na1298_2), .IN3(~na4043_2), .IN4(~na4045_1), .IN5(na1299_1), .IN6(na1300_2),
                      .IN7(na4044_1), .IN8(na1301_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y75     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4043_4 ( .OUT(na4043_2), .IN1(1'b1), .IN2(na1226_2), .IN3(na2992_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x144y79     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4044_1 ( .OUT(na4044_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2984_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na1236_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y82     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4045_1 ( .OUT(na4045_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1227_1), .IN7(na3056_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x142y83     80'h00_0078_00_0000_0CEE_0755
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4054_1 ( .OUT(na4054_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1211_2), .IN6(~na3140_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4054_4 ( .OUT(na4054_2), .IN1(~na1926_1), .IN2(1'b0), .IN3(~na1235_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y79     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4055_1 ( .OUT(na4055_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3048_2), .IN6(1'b1), .IN7(na1222_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x143y84     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4057_4 ( .OUT(na4057_2), .IN1(1'b1), .IN2(na3064_2), .IN3(na1224_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x149y77     80'h00_0018_00_0000_0888_1811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4058_1 ( .OUT(na4058_1), .IN1(~na1309_1), .IN2(~na1306_2), .IN3(~na4061_1), .IN4(~na4059_1), .IN5(na4063_2), .IN6(na4060_1),
                      .IN7(~na4061_2), .IN8(~na4059_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x142y80     80'h00_0078_00_0000_0C88_CA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4059_1 ( .OUT(na4059_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1232_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3073_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4059_4 ( .OUT(na4059_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1208_1), .IN4(na3081_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x145y74     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4060_1 ( .OUT(na4060_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1226_2), .IN7(~na2993_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x140y83     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4061_1 ( .OUT(na4061_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3097_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1230_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4061_4 ( .OUT(na4061_2), .IN1(na2945_1), .IN2(na1229_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x143y79     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4063_4 ( .OUT(na4063_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1235_1), .IN4(~na1927_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x140y72     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4066_1 ( .OUT(na4066_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3141_1), .IN6(1'b1), .IN7(na4260_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x140y77     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4067_4 ( .OUT(na4067_2), .IN1(1'b0), .IN2(~na3009_1), .IN3(~na1220_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x141y77     80'h00_0078_00_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4068_1 ( .OUT(na4068_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3057_1), .IN6(na1227_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4068_4 ( .OUT(na4068_2), .IN1(1'b1), .IN2(na3049_1), .IN3(na1222_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y69     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4071_1 ( .OUT(na4071_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3151_1), .IN8(na1948_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y69     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4072_4 ( .OUT(na4072_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3151_2), .IN4(na1948_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y68     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4073_4 ( .OUT(na4073_2), .IN1(1'b1), .IN2(~na3185_1), .IN3(~na3184_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y71     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4076_4 ( .OUT(na4076_2), .IN1(1'b1), .IN2(~na1334_1), .IN3(na3184_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x88y74     80'h00_0018_00_0000_0CEE_E300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4079_1 ( .OUT(na4079_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3185_1), .IN7(na3184_2), .IN8(na1324_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y78     80'h00_0018_00_0040_0C62_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4082_1 ( .OUT(na4082_1), .IN1(1'b0), .IN2(~na2416_2), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(~na1126_2), .IN7(1'b1), .IN8(na3150_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x131y77     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4083_1 ( .OUT(na4083_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(na1126_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y83     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4085_1 ( .OUT(na4085_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na21_2), .IN6(na57_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y81     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4088_4 ( .OUT(na4088_2), .IN1(1'b1), .IN2(na1126_2), .IN3(1'b1), .IN4(na4196_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y81     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4089_1 ( .OUT(na4089_1), .IN1(1'b1), .IN2(~na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(na4162_2), .IN6(na57_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x129y69     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4093_1 ( .OUT(na4093_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1126_2), .IN7(~na3151_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x109y89     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4100_4 ( .OUT(na4100_2), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(~na24_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x123y65     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4101_1 ( .OUT(na4101_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3131_1), .IN6(~na3133_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y66     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4102_4 ( .OUT(na4102_2), .IN1(na3131_1), .IN2(na3133_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y114     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4103_1 ( .OUT(na4103_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na220_2), .IN6(na221_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y114     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4104_1 ( .OUT(na4104_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na220_2), .IN6(1'b1), .IN7(1'b1), .IN8(na231_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y114     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4105_4 ( .OUT(na4105_2), .IN1(~na226_1), .IN2(1'b1), .IN3(1'b1), .IN4(na230_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y85     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4107_1 ( .OUT(na4107_1), .IN1(1'b1), .IN2(na2416_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2319_1), .IN8(~na2406_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x121y81     80'h00_0060_00_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4109_4 ( .OUT(na4109_2), .IN1(na4107_1), .IN2(~na16_2), .IN3(1'b0), .IN4(na1803_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x108y96     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4110_1 ( .OUT(na4110_1), .IN1(~na1975_2), .IN2(1'b0), .IN3(~na2007_2), .IN4(na19_1), .IN5(~na2039_2), .IN6(~na16_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y82     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4111_4 ( .OUT(na4111_2), .IN1(1'b1), .IN2(~na57_2), .IN3(na215_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y87     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4112_1 ( .OUT(na4112_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4310_2), .IN5(1'b0), .IN6(~na2407_1), .IN7(1'b0), .IN8(~na2320_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x119y85     80'h00_0018_00_0000_0C88_CBFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4114_1 ( .OUT(na4114_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4112_1), .IN6(~na16_2), .IN7(1'b0), .IN8(na1808_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x117y97     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4115_1 ( .OUT(na4115_1), .IN1(~na1976_1), .IN2(1'b0), .IN3(~na2008_1), .IN4(na19_1), .IN5(~na2040_1), .IN6(~na16_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y88     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4116_1 ( .OUT(na4116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na57_2), .IN7(1'b1), .IN8(na263_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y81     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4117_1 ( .OUT(na4117_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na2321_1), .IN7(1'b0), .IN8(~na2408_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x111y79     80'h00_0018_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4119_1 ( .OUT(na4119_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4117_1), .IN6(~na16_2), .IN7(na1813_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x107y90     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4120_1 ( .OUT(na4120_1), .IN1(~na1977_2), .IN2(1'b0), .IN3(~na2009_2), .IN4(na19_1), .IN5(~na2041_2), .IN6(~na16_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y70     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4121_4 ( .OUT(na4121_2), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(na275_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y79     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4122_1 ( .OUT(na4122_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4310_2), .IN5(~na2410_2), .IN6(1'b0), .IN7(~na2323_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x113y79     80'h00_0060_00_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4124_4 ( .OUT(na4124_2), .IN1(na4122_1), .IN2(~na16_2), .IN3(1'b0), .IN4(na1818_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x105y88     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4125_1 ( .OUT(na4125_1), .IN1(~na1979_2), .IN2(1'b0), .IN3(~na2011_2), .IN4(na19_1), .IN5(~na2043_2), .IN6(~na16_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y70     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4126_4 ( .OUT(na4126_2), .IN1(1'b1), .IN2(~na57_2), .IN3(na293_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y83     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4127_1 ( .OUT(na4127_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na2325_1), .IN7(1'b0), .IN8(~na2412_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x111y79     80'h00_0060_00_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4129_4 ( .OUT(na4129_2), .IN1(na4127_1), .IN2(~na16_2), .IN3(1'b0), .IN4(na1823_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x101y88     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4130_1 ( .OUT(na4130_1), .IN1(~na1981_2), .IN2(1'b0), .IN3(~na2013_2), .IN4(na19_1), .IN5(~na2045_2), .IN6(~na16_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y76     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4131_4 ( .OUT(na4131_2), .IN1(na308_1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y79     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4132_1 ( .OUT(na4132_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4310_2), .IN5(1'b0), .IN6(~na2326_2), .IN7(1'b0), .IN8(~na2413_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x117y79     80'h00_0060_00_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4134_4 ( .OUT(na4134_2), .IN1(na4132_1), .IN2(~na16_2), .IN3(1'b0), .IN4(na1828_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x101y78     80'h00_0018_00_0000_0888_F7D3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4135_1 ( .OUT(na4135_1), .IN1(1'b0), .IN2(~na1982_1), .IN3(~na2014_1), .IN4(na19_1), .IN5(~na2046_1), .IN6(~na16_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y74     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4136_1 ( .OUT(na4136_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na312_1), .IN6(~na57_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x144y101     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4141_4 ( .OUT(na4141_2), .IN1(~na3027_1), .IN2(1'b0), .IN3(1'b0), .IN4(na3032_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x147y109     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4146_1 ( .OUT(na4146_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3026_2), .IN8(na891_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x141y117     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4147_1 ( .OUT(na4147_1), .IN1(na963_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na4234_2), .IN6(~na964_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y113     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4151_1 ( .OUT(na4151_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3034_2), .IN6(na964_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y70     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4152_4 ( .OUT(na4152_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na3151_2), .IN4(na1849_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y67     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4153_1 ( .OUT(na4153_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3151_2), .IN8(~na1849_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x160y73     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4154_4 ( .OUT(na4154_2), .IN1(1'b1), .IN2(na3210_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4154_6 ( .RAM_O2(na4154_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4154_2), .COMP_OUT(1'b0) );
// C_///AND/      x107y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4155_4 ( .OUT(na4155_2), .IN1(na1935_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4155_6 ( .RAM_O2(na4155_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4155_2), .COMP_OUT(1'b0) );
// C_///AND/      x111y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4156_4 ( .OUT(na4156_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1934_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4156_6 ( .RAM_O2(na4156_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4156_2), .COMP_OUT(1'b0) );
// C_///AND/      x115y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4157_4 ( .OUT(na4157_2), .IN1(na1935_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4157_6 ( .RAM_O2(na4157_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4157_2), .COMP_OUT(1'b0) );
// C_///AND/      x119y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4158_4 ( .OUT(na4158_2), .IN1(1'b1), .IN2(na1937_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4158_6 ( .RAM_O2(na4158_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4158_2), .COMP_OUT(1'b0) );
// C_///AND/      x123y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4159_4 ( .OUT(na4159_2), .IN1(1'b1), .IN2(na1937_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4159_6 ( .RAM_O2(na4159_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4159_2), .COMP_OUT(1'b0) );
// C_///AND/      x127y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4160_4 ( .OUT(na4160_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1938_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4160_6 ( .RAM_O2(na4160_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4160_2), .COMP_OUT(1'b0) );
// C_////Bridge      x147y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4161_5 ( .OUT(na4161_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4162_5 ( .OUT(na4162_2), .IN1(1'b0), .IN2(na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4163_5 ( .OUT(na4163_2), .IN1(1'b0), .IN2(na16_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y86     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4164_5 ( .OUT(na4164_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y91     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4165_5 ( .OUT(na4165_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na21_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y95     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4166_5 ( .OUT(na4166_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na23_1), .IN8(1'b0) );
// C_////Bridge      x103y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4167_5 ( .OUT(na4167_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na24_2) );
// C_////Bridge      x107y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4168_5 ( .OUT(na4168_2), .IN1(1'b0), .IN2(1'b0), .IN3(na26_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4169_5 ( .OUT(na4169_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4170_5 ( .OUT(na4170_2), .IN1(1'b0), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4171_5 ( .OUT(na4171_2), .IN1(1'b0), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y74     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4172_5 ( .OUT(na4172_2), .IN1(1'b0), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y110     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4173_5 ( .OUT(na4173_2), .IN1(1'b0), .IN2(1'b0), .IN3(na215_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y101     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4174_5 ( .OUT(na4174_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na216_2) );
// C_////Bridge      x122y103     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4175_5 ( .OUT(na4175_2), .IN1(na217_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y112     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4176_5 ( .OUT(na4176_2), .IN1(na219_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y115     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4177_5 ( .OUT(na4177_2), .IN1(1'b0), .IN2(na221_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y114     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4178_5 ( .OUT(na4178_2), .IN1(1'b0), .IN2(na221_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y106     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4179_5 ( .OUT(na4179_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na222_2), .IN8(1'b0) );
// C_////Bridge      x123y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4180_5 ( .OUT(na4180_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na227_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x130y112     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4181_5 ( .OUT(na4181_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na232_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y110     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4182_5 ( .OUT(na4182_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na239_1) );
// C_////Bridge      x124y110     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4183_5 ( .OUT(na4183_2), .IN1(1'b0), .IN2(1'b0), .IN3(na242_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y112     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4184_5 ( .OUT(na4184_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na244_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y108     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4185_5 ( .OUT(na4185_2), .IN1(1'b0), .IN2(na245_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y106     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4186_5 ( .OUT(na4186_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na247_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y110     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4187_5 ( .OUT(na4187_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na248_1) );
// C_////Bridge      x121y112     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4188_5 ( .OUT(na4188_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na269_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y111     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4189_5 ( .OUT(na4189_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na270_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4190_5 ( .OUT(na4190_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na275_1) );
// C_////Bridge      x106y78     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4191_5 ( .OUT(na4191_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na294_1), .IN8(1'b0) );
// C_////Bridge      x138y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4192_5 ( .OUT(na4192_2), .IN1(1'b0), .IN2(1'b0), .IN3(na322_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x141y68     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4193_5 ( .OUT(na4193_2), .IN1(1'b0), .IN2(1'b0), .IN3(na322_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4194_5 ( .OUT(na4194_2), .IN1(na323_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4195_5 ( .OUT(na4195_2), .IN1(na323_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y80     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4196_5 ( .OUT(na4196_2), .IN1(1'b0), .IN2(na543_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y114     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4197_5 ( .OUT(na4197_2), .IN1(1'b0), .IN2(1'b0), .IN3(na800_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x146y112     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4198_5 ( .OUT(na4198_2), .IN1(na811_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y114     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4199_5 ( .OUT(na4199_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na812_2), .IN8(1'b0) );
// C_////Bridge      x151y113     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4200_5 ( .OUT(na4200_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na813_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x152y113     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4201_5 ( .OUT(na4201_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na814_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y113     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4202_5 ( .OUT(na4202_2), .IN1(1'b0), .IN2(1'b0), .IN3(na815_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y115     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4203_5 ( .OUT(na4203_2), .IN1(1'b0), .IN2(na816_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y110     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4204_5 ( .OUT(na4204_2), .IN1(1'b0), .IN2(na818_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y116     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4205_5 ( .OUT(na4205_2), .IN1(1'b0), .IN2(na819_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y108     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4206_5 ( .OUT(na4206_2), .IN1(na823_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y107     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4207_5 ( .OUT(na4207_2), .IN1(1'b0), .IN2(1'b0), .IN3(na832_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y106     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4208_5 ( .OUT(na4208_2), .IN1(1'b0), .IN2(na833_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y107     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4209_5 ( .OUT(na4209_2), .IN1(1'b0), .IN2(1'b0), .IN3(na836_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y112     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4210_5 ( .OUT(na4210_2), .IN1(na843_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y108     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4211_5 ( .OUT(na4211_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na847_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y105     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4212_5 ( .OUT(na4212_2), .IN1(1'b0), .IN2(na855_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x130y74     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4213_5 ( .OUT(na4213_2), .IN1(1'b0), .IN2(na856_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y114     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4214_5 ( .OUT(na4214_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na864_1) );
// C_////Bridge      x108y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4215_5 ( .OUT(na4215_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na875_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y107     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4216_5 ( .OUT(na4216_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na879_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y99     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4217_5 ( .OUT(na4217_2), .IN1(1'b0), .IN2(1'b0), .IN3(na888_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4218_5 ( .OUT(na4218_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na891_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4219_5 ( .OUT(na4219_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na893_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y109     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4220_5 ( .OUT(na4220_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na893_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x151y112     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4221_5 ( .OUT(na4221_2), .IN1(1'b0), .IN2(1'b0), .IN3(na900_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y100     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4222_5 ( .OUT(na4222_2), .IN1(na903_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y94     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4223_5 ( .OUT(na4223_2), .IN1(na903_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y97     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4224_5 ( .OUT(na4224_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na906_1) );
// C_////Bridge      x147y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4225_5 ( .OUT(na4225_2), .IN1(na908_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y103     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4226_5 ( .OUT(na4226_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na911_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y101     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4227_5 ( .OUT(na4227_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na919_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4228_5 ( .OUT(na4228_2), .IN1(1'b0), .IN2(na924_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x142y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4229_5 ( .OUT(na4229_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4230_5 ( .OUT(na4230_2), .IN1(1'b0), .IN2(na933_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y83     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4231_5 ( .OUT(na4231_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na949_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y116     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4232_5 ( .OUT(na4232_2), .IN1(na963_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x131y115     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4233_5 ( .OUT(na4233_2), .IN1(1'b0), .IN2(na964_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y117     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4234_5 ( .OUT(na4234_2), .IN1(1'b0), .IN2(1'b0), .IN3(na965_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y116     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4235_5 ( .OUT(na4235_2), .IN1(1'b0), .IN2(1'b0), .IN3(na965_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y117     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4236_5 ( .OUT(na4236_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na967_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4237_5 ( .OUT(na4237_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na969_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y118     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4238_5 ( .OUT(na4238_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na970_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y112     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4239_5 ( .OUT(na4239_2), .IN1(1'b0), .IN2(na974_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x133y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4240_5 ( .OUT(na4240_2), .IN1(na975_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y115     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4241_5 ( .OUT(na4241_2), .IN1(na975_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x131y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4242_5 ( .OUT(na4242_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na983_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y112     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4243_5 ( .OUT(na4243_2), .IN1(1'b0), .IN2(na984_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x129y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4244_5 ( .OUT(na4244_2), .IN1(na988_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y117     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4245_5 ( .OUT(na4245_2), .IN1(na988_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4246_5 ( .OUT(na4246_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na996_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y111     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4247_5 ( .OUT(na4247_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na996_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4248_5 ( .OUT(na4248_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na996_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x135y108     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4249_5 ( .OUT(na4249_2), .IN1(na998_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y108     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4250_5 ( .OUT(na4250_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1001_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y109     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4251_5 ( .OUT(na4251_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1003_1) );
// C_////Bridge      x120y110     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4252_5 ( .OUT(na4252_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1005_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y100     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4253_5 ( .OUT(na4253_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1014_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4254_5 ( .OUT(na4254_2), .IN1(na1026_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x135y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4255_5 ( .OUT(na4255_2), .IN1(1'b0), .IN2(na1126_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4256_5 ( .OUT(na4256_2), .IN1(1'b0), .IN2(na1126_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4257_5 ( .OUT(na4257_2), .IN1(1'b0), .IN2(na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4258_5 ( .OUT(na4258_2), .IN1(1'b0), .IN2(na1136_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4259_5 ( .OUT(na4259_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1206_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4260_5 ( .OUT(na4260_2), .IN1(na1211_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y79     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4261_5 ( .OUT(na4261_2), .IN1(na1219_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4262_5 ( .OUT(na4262_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1220_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4263_5 ( .OUT(na4263_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1222_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x142y90     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4264_5 ( .OUT(na4264_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1224_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4265_5 ( .OUT(na4265_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1232_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y78     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4266_5 ( .OUT(na4266_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1233_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4267_5 ( .OUT(na4267_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1236_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4268_5 ( .OUT(na4268_2), .IN1(na1319_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4269_5 ( .OUT(na4269_2), .IN1(na1319_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4270_5 ( .OUT(na4270_2), .IN1(1'b0), .IN2(na1325_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y64     80'h00_00A2_24_7000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4271_5 ( .OUT(na4271_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1357_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4272_5 ( .OUT(na4272_2), .IN1(na1358_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4273_5 ( .OUT(na4273_2), .IN1(1'b0), .IN2(na1376_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4274_5 ( .OUT(na4274_2), .IN1(1'b0), .IN2(na1376_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4275_5 ( .OUT(na4275_2), .IN1(1'b0), .IN2(na1387_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4276_5 ( .OUT(na4276_2), .IN1(1'b0), .IN2(na1387_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4277_5 ( .OUT(na4277_2), .IN1(1'b0), .IN2(na1406_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4278_5 ( .OUT(na4278_2), .IN1(1'b0), .IN2(na1406_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y68     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4279_5 ( .OUT(na4279_2), .IN1(1'b0), .IN2(na1468_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y113     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4280_5 ( .OUT(na4280_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1483_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y103     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4281_5 ( .OUT(na4281_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1490_2) );
// C_////Bridge      x134y114     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4282_5 ( .OUT(na4282_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1799_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y113     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4283_5 ( .OUT(na4283_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1801_1) );
// C_////Bridge      x145y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4284_5 ( .OUT(na4284_2), .IN1(na1834_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4285_5 ( .OUT(na4285_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1836_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x142y111     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4286_5 ( .OUT(na4286_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1836_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y104     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4287_5 ( .OUT(na4287_2), .IN1(na1839_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x146y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4288_5 ( .OUT(na4288_2), .IN1(na1839_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y102     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4289_5 ( .OUT(na4289_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1841_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y103     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4290_5 ( .OUT(na4290_2), .IN1(1'b0), .IN2(na1843_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x133y116     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4291_5 ( .OUT(na4291_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1846_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y116     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4292_5 ( .OUT(na4292_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1846_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4293_5 ( .OUT(na4293_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1848_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x133y118     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4294_5 ( .OUT(na4294_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1848_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4295_5 ( .OUT(na4295_2), .IN1(1'b0), .IN2(na1922_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y69     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4296_5 ( .OUT(na4296_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1930_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y96     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4297_5 ( .OUT(na4297_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1935_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y95     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4298_5 ( .OUT(na4298_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1935_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4299_5 ( .OUT(na4299_2), .IN1(1'b0), .IN2(na1937_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4300_5 ( .OUT(na4300_2), .IN1(1'b0), .IN2(na1941_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y94     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4301_5 ( .OUT(na4301_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1943_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4302_5 ( .OUT(na4302_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1947_2), .IN8(1'b0) );
// C_////Bridge      x132y68     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4303_5 ( .OUT(na4303_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1957_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y87     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4304_5 ( .OUT(na4304_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1958_1), .IN8(1'b0) );
// C_////Bridge      x88y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4305_5 ( .OUT(na4305_2), .IN1(na2283_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y108     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4306_5 ( .OUT(na4306_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2287_1), .IN8(1'b0) );
// C_////Bridge      x110y80     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4307_5 ( .OUT(na4307_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2292_2), .IN8(1'b0) );
// C_////Bridge      x131y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4308_5 ( .OUT(na4308_2), .IN1(1'b0), .IN2(na2296_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4309_5 ( .OUT(na4309_2), .IN1(na2415_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y88     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4310_5 ( .OUT(na4310_2), .IN1(1'b0), .IN2(na2416_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4311_5 ( .OUT(na4311_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2418_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y98     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4312_5 ( .OUT(na4312_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2419_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4313_5 ( .OUT(na4313_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2419_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y100     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4314_5 ( .OUT(na4314_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2421_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4315_5 ( .OUT(na4315_2), .IN1(1'b0), .IN2(na2422_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4316_5 ( .OUT(na4316_2), .IN1(1'b0), .IN2(na2423_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y77     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4317_5 ( .OUT(na4317_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2433_2), .IN8(1'b0) );
// C_////Bridge      x119y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4318_5 ( .OUT(na4318_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2438_1) );
// C_////Bridge      x88y93     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4319_5 ( .OUT(na4319_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2447_1) );
// C_////Bridge      x109y90     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4320_5 ( .OUT(na4320_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2449_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4321_5 ( .OUT(na4321_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2449_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y98     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4322_5 ( .OUT(na4322_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2453_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4323_5 ( .OUT(na4323_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2453_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y92     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4324_5 ( .OUT(na4324_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2456_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y94     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4325_5 ( .OUT(na4325_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2457_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y83     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4326_5 ( .OUT(na4326_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2460_2), .IN8(1'b0) );
// C_////Bridge      x118y83     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4327_5 ( .OUT(na4327_2), .IN1(na2463_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y64     80'h00_00A6_24_7000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4328_5 ( .OUT(na4328_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2465_2), .IN8(1'b0) );
// C_////Bridge      x128y96     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4329_5 ( .OUT(na4329_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2467_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y97     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4330_5 ( .OUT(na4330_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2468_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4331_5 ( .OUT(na4331_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2470_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y93     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4332_5 ( .OUT(na4332_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2472_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x133y100     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4333_5 ( .OUT(na4333_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2475_1), .IN8(1'b0) );
// C_////Bridge      x119y110     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4334_5 ( .OUT(na4334_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2477_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y86     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4335_5 ( .OUT(na4335_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2761_1), .IN8(1'b0) );
// C_////Bridge      x100y101     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4336_5 ( .OUT(na4336_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2770_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4337_5 ( .OUT(na4337_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2774_2) );
// C_////Bridge      x110y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4338_5 ( .OUT(na4338_2), .IN1(1'b0), .IN2(na2784_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y83     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4339_5 ( .OUT(na4339_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2793_1) );
// C_////Bridge      x107y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4340_5 ( .OUT(na4340_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2797_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y96     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4341_5 ( .OUT(na4341_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2801_1), .IN8(1'b0) );
// C_////Bridge      x129y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4342_5 ( .OUT(na4342_2), .IN1(na2846_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y113     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4343_5 ( .OUT(na4343_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2867_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y114     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4344_5 ( .OUT(na4344_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2892_2), .IN8(1'b0) );
// C_////Bridge      x94y92     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4345_5 ( .OUT(na4345_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2895_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4346_5 ( .OUT(na4346_2), .IN1(na2905_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4347_5 ( .OUT(na4347_2), .IN1(1'b0), .IN2(na2946_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y69     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4348_5 ( .OUT(na4348_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2956_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4349_5 ( .OUT(na4349_2), .IN1(na2961_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4350_5 ( .OUT(na4350_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2967_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y68     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4351_5 ( .OUT(na4351_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2969_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4352_5 ( .OUT(na4352_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2970_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4353_5 ( .OUT(na4353_2), .IN1(na2985_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4354_5 ( .OUT(na4354_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3000_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y107     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4355_5 ( .OUT(na4355_2), .IN1(na3010_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4356_5 ( .OUT(na4356_2), .IN1(na3010_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x133y110     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4357_5 ( .OUT(na4357_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3011_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x132y110     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4358_5 ( .OUT(na4358_2), .IN1(na3017_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y115     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4359_5 ( .OUT(na4359_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3018_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y112     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4360_5 ( .OUT(na4360_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3019_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y114     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4361_5 ( .OUT(na4361_2), .IN1(1'b0), .IN2(na3022_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y112     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4362_5 ( .OUT(na4362_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3023_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y112     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4363_5 ( .OUT(na4363_2), .IN1(na3025_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y110     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4364_5 ( .OUT(na4364_2), .IN1(na3025_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y110     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4365_5 ( .OUT(na4365_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3026_2), .IN8(1'b0) );
// C_////Bridge      x150y97     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4366_5 ( .OUT(na4366_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3027_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y101     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4367_5 ( .OUT(na4367_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3031_2) );
// C_////Bridge      x149y98     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4368_5 ( .OUT(na4368_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3032_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4369_5 ( .OUT(na4369_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3033_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y102     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4370_5 ( .OUT(na4370_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3033_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y100     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4371_5 ( .OUT(na4371_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3033_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4372_5 ( .OUT(na4372_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3033_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y111     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4373_5 ( .OUT(na4373_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3035_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y115     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4374_5 ( .OUT(na4374_2), .IN1(1'b0), .IN2(na3038_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y114     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4375_5 ( .OUT(na4375_2), .IN1(1'b0), .IN2(na3038_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y113     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4376_5 ( .OUT(na4376_2), .IN1(na3039_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4377_5 ( .OUT(na4377_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3041_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4378_5 ( .OUT(na4378_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3041_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4379_5 ( .OUT(na4379_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3137_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y79     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4380_5 ( .OUT(na4380_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3150_2) );
// C_////Bridge      x131y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4381_5 ( .OUT(na4381_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3151_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4382_5 ( .OUT(na4382_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3151_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x132y64     80'h00_00A2_24_7000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4383_5 ( .OUT(na4383_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3151_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4384_5 ( .OUT(na4384_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3170_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y69     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4385_5 ( .OUT(na4385_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3170_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y69     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4386_5 ( .OUT(na4386_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3174_2), .IN8(1'b0) );
// C_////Bridge      x92y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4387_5 ( .OUT(na4387_2), .IN1(1'b0), .IN2(na3181_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y79     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4388_5 ( .OUT(na4388_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3184_2), .IN8(1'b0) );
// C_////Bridge      x93y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4389_5 ( .OUT(na4389_2), .IN1(1'b0), .IN2(na3185_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4390_5 ( .OUT(na4390_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3211_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4391_5 ( .OUT(na4391_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3223_1), .IN8(1'b0) );
// C_////Bridge      x145y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4392_5 ( .OUT(na4392_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3223_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x142y74     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4393_5 ( .OUT(na4393_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3234_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4394_5 ( .OUT(na4394_2), .IN1(na3235_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y98     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4395_5 ( .OUT(na4395_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3278_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y109     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4396_5 ( .OUT(na4396_2), .IN1(na3442_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x131y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4397_5 ( .OUT(na4397_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3570_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y85     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4398_5 ( .OUT(na4398_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3663_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y116     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4399_5 ( .OUT(na4399_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3700_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4400_5 ( .OUT(na4400_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3704_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x142y113     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4401_5 ( .OUT(na4401_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3709_1) );
// C_////Bridge      x147y108     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4402_5 ( .OUT(na4402_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3712_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y99     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4403_5 ( .OUT(na4403_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3739_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y113     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4404_5 ( .OUT(na4404_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3781_1) );
// C_////Bridge      x135y115     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4405_5 ( .OUT(na4405_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3790_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x131y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4406_5 ( .OUT(na4406_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3796_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4407_5 ( .OUT(na4407_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3863_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y94     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4408_5 ( .OUT(na4408_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3864_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y80     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4409_5 ( .OUT(na4409_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3865_2), .IN8(1'b0) );
// C_////Bridge      x122y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4410_5 ( .OUT(na4410_2), .IN1(na3866_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y74     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4411_5 ( .OUT(na4411_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3867_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4412_5 ( .OUT(na4412_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3868_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4413_5 ( .OUT(na4413_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3869_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y79     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4414_5 ( .OUT(na4414_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3870_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4415_5 ( .OUT(na4415_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4068_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x130y64     80'h00_00A0_24_7000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4416_5 ( .OUT(na4416_2), .IN1(na4153_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_CP_route////      x83y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4417_1 ( .OUT(na4417_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x84y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4418_1 ( .OUT(na4418_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x85y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4419_1 ( .OUT(na4419_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x86y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4420_1 ( .OUT(na4420_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x87y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4421_1 ( .OUT(na4421_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x88y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4422_1 ( .OUT(na4422_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x89y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4423_1 ( .OUT(na4423_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x90y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4424_1 ( .OUT(na4424_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x91y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4425_1 ( .OUT(na4425_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x92y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4426_1 ( .OUT(na4426_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x93y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4427_1 ( .OUT(na4427_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x95y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4428_1 ( .OUT(na4428_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x96y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4429_1 ( .OUT(na4429_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x97y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4430_1 ( .OUT(na4430_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x98y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4431_1 ( .OUT(na4431_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x99y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4432_1 ( .OUT(na4432_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x100y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4433_1 ( .OUT(na4433_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x101y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4434_1 ( .OUT(na4434_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x102y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4435_1 ( .OUT(na4435_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x103y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4436_1 ( .OUT(na4436_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x104y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4437_1 ( .OUT(na4437_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x105y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4438_1 ( .OUT(na4438_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x106y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4439_1 ( .OUT(na4439_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x107y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4440_1 ( .OUT(na4440_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x108y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4441_1 ( .OUT(na4441_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x109y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4442_1 ( .OUT(na4442_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x110y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4443_1 ( .OUT(na4443_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x111y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4444_1 ( .OUT(na4444_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x112y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4445_1 ( .OUT(na4445_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x113y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4446_1 ( .OUT(na4446_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x114y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4447_1 ( .OUT(na4447_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x115y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4448_1 ( .OUT(na4448_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x116y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4449_1 ( .OUT(na4449_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x117y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4450_1 ( .OUT(na4450_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x118y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4451_1 ( .OUT(na4451_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x119y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4452_1 ( .OUT(na4452_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x120y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4453_1 ( .OUT(na4453_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x121y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4454_1 ( .OUT(na4454_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x122y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4455_1 ( .OUT(na4455_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x123y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4456_1 ( .OUT(na4456_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x124y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4457_1 ( .OUT(na4457_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x125y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4458_1 ( .OUT(na4458_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x126y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4459_1 ( .OUT(na4459_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x127y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4460_1 ( .OUT(na4460_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x128y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4461_1 ( .OUT(na4461_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x129y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4462_1 ( .OUT(na4462_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x131y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4463_1 ( .OUT(na4463_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x133y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4464_1 ( .OUT(na4464_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x134y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4465_1 ( .OUT(na4465_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x135y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4466_1 ( .OUT(na4466_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x136y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4467_1 ( .OUT(na4467_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x137y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4468_1 ( .OUT(na4468_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x138y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4469_1 ( .OUT(na4469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x139y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4470_1 ( .OUT(na4470_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x140y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4471_1 ( .OUT(na4471_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x141y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4472_1 ( .OUT(na4472_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x142y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4473_1 ( .OUT(na4473_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x143y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4474_1 ( .OUT(na4474_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x144y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4475_1 ( .OUT(na4475_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x145y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4476_1 ( .OUT(na4476_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x146y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4477_1 ( .OUT(na4477_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x147y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4478_1 ( .OUT(na4478_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x149y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4479_1 ( .OUT(na4479_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x150y64     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4480_1 ( .OUT(na4480_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x82y64     80'h00_0078_09_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4481_1 ( .OUT(na4481_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1928_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4481_4 ( .OUT(na4481_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9000)) 
           _a4481_6 ( .COUTX(na4481_3), .POUTX(na4481_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na4481_1), .OUT2(na4481_2), .COMP_OUT(1'b0) );
endmodule
