//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 Jul 2023)
//  Compile Time: 2023-07-20 13:23:25
//  Program Run:  2023-08-07 04:10:11
//  Program Call: ../../bin/p_r/p_r -i net/aes256_uart_synth.v -o aes256_uart -ccf src/aes256_uart.ccf 
//  File Type:    Verilog

// Gatecount:   2872
module aes256_uart (clk , data_in , reset_n ,
       data_out , led 
       ) ;

input  clk;
input  data_in;
input  reset_n;

output data_out;
output [5:0]led;



wire [5:0]led;
wire clk;
wire data_in;
wire na1_1;
wire na2_1;
wire na2_1_i;
wire na3_1;
wire na3_1_i;
wire na3_2;
wire na3_2_i;
wire na5_1;
wire na5_1_i;
wire na5_2;
wire na5_2_i;
wire na6_1;
wire na6_1_i;
wire na7_1;
wire na9_2;
wire na9_2_i;
wire na10_1;
wire na10_1_i;
wire na10_2;
wire na10_2_i;
wire na12_1;
wire na12_1_i;
wire na12_2;
wire na12_2_i;
wire na13_1;
wire na13_1_i;
wire na14_1;
wire na15_2;
wire na16_2;
wire na17_1;
wire na21_1;
wire na21_2;
wire na22_1;
wire na24_1;
wire na25_1;
wire na25_2;
wire na26_1;
wire na26_2;
wire na27_1;
wire na27_1_i;
wire na28_1;
wire na30_1;
wire na32_1;
wire na33_1;
wire na34_1;
wire na34_1_i;
wire na35_2;
wire na36_1;
wire na38_1;
wire na39_1;
wire na40_1;
wire na40_1_i;
wire na41_1;
wire na42_1;
wire na44_1;
wire na45_1;
wire na46_1;
wire na46_1_i;
wire na47_2;
wire na48_1;
wire na50_1;
wire na51_1;
wire na52_1;
wire na52_1_i;
wire na53_1;
wire na54_1;
wire na56_1;
wire na57_1;
wire na58_1;
wire na58_1_i;
wire na59_2;
wire na60_1;
wire na62_1;
wire na63_1;
wire na64_1;
wire na64_1_i;
wire na65_1;
wire na66_1;
wire na68_1;
wire na69_1;
wire na70_1;
wire na70_1_i;
wire na71_2;
wire na72_1;
wire na74_1;
wire na75_1;
wire na76_1;
wire na76_1_i;
wire na77_1;
wire na78_1;
wire na80_1;
wire na81_1;
wire na82_1;
wire na82_1_i;
wire na83_2;
wire na84_1;
wire na86_1;
wire na87_1;
wire na88_1;
wire na88_1_i;
wire na89_1;
wire na90_1;
wire na92_1;
wire na93_1;
wire na94_1;
wire na94_1_i;
wire na95_2;
wire na96_1;
wire na98_1;
wire na99_1;
wire na100_1;
wire na100_1_i;
wire na101_1;
wire na102_1;
wire na104_1;
wire na105_1;
wire na106_1;
wire na106_1_i;
wire na107_2;
wire na108_1;
wire na110_1;
wire na111_1;
wire na112_1;
wire na112_1_i;
wire na113_1;
wire na114_1;
wire na116_1;
wire na117_1;
wire na118_1;
wire na118_1_i;
wire na119_2;
wire na120_1;
wire na122_1;
wire na123_1;
wire na124_1;
wire na124_1_i;
wire na125_1;
wire na126_1;
wire na128_1;
wire na129_1;
wire na130_1;
wire na130_1_i;
wire na131_2;
wire na132_1;
wire na134_1;
wire na135_1;
wire na136_1;
wire na136_1_i;
wire na137_1;
wire na138_1;
wire na140_1;
wire na141_1;
wire na142_1;
wire na142_1_i;
wire na143_2;
wire na144_1;
wire na146_1;
wire na147_1;
wire na148_1;
wire na148_1_i;
wire na149_1;
wire na150_1;
wire na152_1;
wire na153_1;
wire na154_1;
wire na154_1_i;
wire na155_2;
wire na156_1;
wire na158_1;
wire na159_1;
wire na160_1;
wire na160_1_i;
wire na161_1;
wire na162_1;
wire na164_1;
wire na165_1;
wire na166_1;
wire na166_1_i;
wire na167_2;
wire na168_1;
wire na170_1;
wire na171_1;
wire na172_1;
wire na172_1_i;
wire na173_1;
wire na174_1;
wire na176_1;
wire na177_1;
wire na178_1;
wire na178_1_i;
wire na179_2;
wire na180_1;
wire na182_1;
wire na183_1;
wire na184_1;
wire na184_1_i;
wire na185_1;
wire na186_1;
wire na188_1;
wire na189_1;
wire na190_1;
wire na190_1_i;
wire na191_2;
wire na192_1;
wire na194_1;
wire na195_1;
wire na196_1;
wire na196_1_i;
wire na197_1;
wire na198_1;
wire na200_1;
wire na201_1;
wire na202_1;
wire na202_1_i;
wire na203_2;
wire na204_1;
wire na206_1;
wire na207_1;
wire na208_1;
wire na208_1_i;
wire na209_1;
wire na210_1;
wire na212_1;
wire na213_1;
wire na214_1;
wire na214_2;
wire na215_1;
wire na215_2;
wire na216_1;
wire na217_1;
wire na218_1;
wire na221_1;
wire na223_2;
wire na225_1;
wire na225_2;
wire na227_1;
wire na228_1;
wire na229_1;
wire na231_1;
wire na233_2;
wire na234_1;
wire na236_1;
wire na238_1;
wire na239_1;
wire na240_2;
wire na241_1;
wire na242_2;
wire na243_1;
wire na244_1;
wire na245_1;
wire na246_1;
wire na248_2;
wire na249_2;
wire na250_1;
wire na251_1;
wire na252_1;
wire na253_1;
wire na254_1;
wire na255_1;
wire na256_1;
wire na259_1;
wire na260_1;
wire na261_2;
wire na262_1;
wire na263_1;
wire na264_1;
wire na264_2;
wire na265_1;
wire na267_1;
wire na268_1;
wire na269_1;
wire na271_1;
wire na272_1;
wire na273_1;
wire na274_1;
wire na275_1;
wire na276_2;
wire na277_1;
wire na277_2;
wire na278_1;
wire na279_1;
wire na279_1_i;
wire na280_1;
wire na282_1;
wire na283_1;
wire na284_1;
wire na285_1;
wire na287_1;
wire na287_2;
wire na290_1;
wire na291_1;
wire na292_2;
wire na293_1;
wire na294_2;
wire na295_1;
wire na295_2;
wire na296_1;
wire na297_1;
wire na298_1;
wire na299_2;
wire na300_1;
wire na300_2;
wire na301_2;
wire na303_2;
wire na304_1;
wire na306_1;
wire na307_1;
wire na308_1;
wire na309_1;
wire na309_2;
wire na310_1;
wire na311_1;
wire na312_1;
wire na313_1;
wire na314_2;
wire na315_1;
wire na315_2;
wire na316_1;
wire na316_1_i;
wire na317_1;
wire na319_1;
wire na320_1;
wire na321_1;
wire na322_1;
wire na324_1;
wire na324_1_i;
wire na325_1;
wire na327_1;
wire na328_1;
wire na329_1;
wire na330_1;
wire na333_1;
wire na333_1_i;
wire na334_1;
wire na336_1;
wire na337_1;
wire na338_1;
wire na339_1;
wire na342_1;
wire na342_1_i;
wire na343_1;
wire na345_1;
wire na346_1;
wire na349_1;
wire na349_2;
wire na350_1;
wire na353_1;
wire na353_1_i;
wire na354_1;
wire na356_1;
wire na357_1;
wire na359_1;
wire na362_1;
wire na362_1_i;
wire na363_1;
wire na365_1;
wire na366_1;
wire na367_1;
wire na368_1;
wire na371_1;
wire na371_1_i;
wire na374_1;
wire na378_1;
wire na379_1;
wire na380_1;
wire na380_1_i;
wire na381_1;
wire na383_1;
wire na384_1;
wire na386_1;
wire na389_1;
wire na389_1_i;
wire na390_1;
wire na392_1;
wire na393_1;
wire na397_1;
wire na397_1_i;
wire na398_1;
wire na400_1;
wire na401_1;
wire na405_1;
wire na405_1_i;
wire na406_1;
wire na408_1;
wire na409_1;
wire na410_1;
wire na411_1;
wire na414_1;
wire na414_1_i;
wire na415_1;
wire na417_1;
wire na418_1;
wire na420_1;
wire na423_1;
wire na423_1_i;
wire na426_1;
wire na430_1;
wire na431_1;
wire na432_1;
wire na432_1_i;
wire na433_1;
wire na437_1;
wire na439_1;
wire na440_1;
wire na441_1;
wire na441_1_i;
wire na442_1;
wire na444_1;
wire na445_1;
wire na449_1;
wire na449_1_i;
wire na450_1;
wire na452_1;
wire na453_1;
wire na455_1;
wire na458_1;
wire na458_1_i;
wire na461_1;
wire na465_1;
wire na466_1;
wire na467_1;
wire na467_1_i;
wire na468_1;
wire na470_1;
wire na471_1;
wire na472_1;
wire na473_1;
wire na476_1;
wire na476_1_i;
wire na477_1;
wire na481_2;
wire na483_1;
wire na484_1;
wire na485_1;
wire na485_1_i;
wire na486_1;
wire na488_1;
wire na489_1;
wire na491_1;
wire na494_1;
wire na494_1_i;
wire na495_1;
wire na497_1;
wire na498_1;
wire na500_1;
wire na503_1;
wire na503_1_i;
wire na504_1;
wire na506_1;
wire na507_1;
wire na508_2;
wire na509_1;
wire na512_1;
wire na512_1_i;
wire na515_1;
wire na519_1;
wire na520_1;
wire na521_1;
wire na521_1_i;
wire na522_1;
wire na524_1;
wire na525_1;
wire na527_1;
wire na530_1;
wire na530_1_i;
wire na531_1;
wire na533_1;
wire na534_1;
wire na535_1;
wire na536_1;
wire na539_1;
wire na539_1_i;
wire na540_1;
wire na541_1;
wire na542_2;
wire na543_2;
wire na544_1;
wire na545_2;
wire na546_2;
wire na547_1;
wire na548_2;
wire na548_2_i;
wire na549_1;
wire na549_1_i;
wire na550_1;
wire na551_1;
wire na551_1_i;
wire na552_2;
wire na553_1;
wire na553_1_i;
wire na554_1;
wire na554_1_i;
wire na555_1;
wire na555_1_i;
wire na556_1;
wire na556_1_i;
wire na557_1;
wire na557_1_i;
wire na558_1;
wire na558_1_i;
wire na559_1;
wire na559_1_i;
wire na560_1;
wire na560_1_i;
wire na561_1;
wire na561_1_i;
wire na562_1;
wire na562_1_i;
wire na563_1;
wire na563_1_i;
wire na564_1;
wire na564_1_i;
wire na565_1;
wire na565_1_i;
wire na566_1;
wire na566_1_i;
wire na567_1;
wire na567_1_i;
wire na568_1;
wire na568_1_i;
wire na569_1;
wire na569_1_i;
wire na570_1;
wire na570_1_i;
wire na571_1;
wire na571_1_i;
wire na572_1;
wire na572_1_i;
wire na573_1;
wire na573_1_i;
wire na574_1;
wire na574_1_i;
wire na575_1;
wire na575_1_i;
wire na576_1;
wire na576_1_i;
wire na577_1;
wire na577_1_i;
wire na578_1;
wire na578_1_i;
wire na579_1;
wire na579_1_i;
wire na580_1;
wire na580_1_i;
wire na581_1;
wire na581_1_i;
wire na582_1;
wire na582_1_i;
wire na583_1;
wire na583_1_i;
wire na584_1;
wire na584_1_i;
wire na585_1;
wire na585_1_i;
wire na586_1;
wire na586_1_i;
wire na587_1;
wire na587_1_i;
wire na588_1;
wire na588_1_i;
wire na589_1;
wire na589_1_i;
wire na590_1;
wire na590_1_i;
wire na591_1;
wire na591_1_i;
wire na592_1;
wire na592_1_i;
wire na593_1;
wire na593_1_i;
wire na594_1;
wire na594_1_i;
wire na595_1;
wire na595_1_i;
wire na596_1;
wire na596_1_i;
wire na597_1;
wire na597_1_i;
wire na598_1;
wire na598_1_i;
wire na599_1;
wire na599_1_i;
wire na600_1;
wire na600_1_i;
wire na601_1;
wire na601_1_i;
wire na602_1;
wire na602_1_i;
wire na603_1;
wire na603_1_i;
wire na604_1;
wire na604_1_i;
wire na605_1;
wire na605_1_i;
wire na606_1;
wire na606_1_i;
wire na607_1;
wire na607_1_i;
wire na608_1;
wire na608_1_i;
wire na609_1;
wire na609_1_i;
wire na610_1;
wire na610_1_i;
wire na611_1;
wire na611_1_i;
wire na612_1;
wire na612_1_i;
wire na613_1;
wire na613_1_i;
wire na614_1;
wire na614_1_i;
wire na615_1;
wire na615_1_i;
wire na616_1;
wire na616_1_i;
wire na617_1;
wire na617_1_i;
wire na618_1;
wire na618_1_i;
wire na619_1;
wire na619_1_i;
wire na620_1;
wire na620_1_i;
wire na621_1;
wire na621_1_i;
wire na622_1;
wire na622_1_i;
wire na623_1;
wire na623_1_i;
wire na624_1;
wire na624_1_i;
wire na625_1;
wire na625_1_i;
wire na626_1;
wire na626_1_i;
wire na627_1;
wire na627_1_i;
wire na628_1;
wire na628_1_i;
wire na629_1;
wire na629_1_i;
wire na630_1;
wire na630_1_i;
wire na631_1;
wire na631_1_i;
wire na632_1;
wire na632_1_i;
wire na633_1;
wire na633_1_i;
wire na634_1;
wire na634_1_i;
wire na635_1;
wire na635_1_i;
wire na636_1;
wire na636_1_i;
wire na637_1;
wire na637_1_i;
wire na638_1;
wire na638_1_i;
wire na639_1;
wire na639_1_i;
wire na640_1;
wire na640_1_i;
wire na641_1;
wire na641_1_i;
wire na642_1;
wire na642_1_i;
wire na643_1;
wire na643_1_i;
wire na644_1;
wire na644_1_i;
wire na645_1;
wire na645_1_i;
wire na646_1;
wire na646_1_i;
wire na647_1;
wire na647_1_i;
wire na648_1;
wire na648_1_i;
wire na649_1;
wire na649_1_i;
wire na650_1;
wire na650_1_i;
wire na651_1;
wire na651_1_i;
wire na652_1;
wire na652_1_i;
wire na653_1;
wire na653_1_i;
wire na654_1;
wire na654_1_i;
wire na655_1;
wire na655_1_i;
wire na656_1;
wire na656_1_i;
wire na657_1;
wire na657_1_i;
wire na658_1;
wire na658_1_i;
wire na659_1;
wire na659_1_i;
wire na660_1;
wire na660_1_i;
wire na661_1;
wire na661_1_i;
wire na662_1;
wire na662_1_i;
wire na663_1;
wire na663_1_i;
wire na664_1;
wire na664_1_i;
wire na665_1;
wire na665_1_i;
wire na666_1;
wire na666_1_i;
wire na667_1;
wire na667_1_i;
wire na668_1;
wire na668_1_i;
wire na669_1;
wire na669_1_i;
wire na670_1;
wire na670_1_i;
wire na671_1;
wire na671_1_i;
wire na672_1;
wire na672_1_i;
wire na673_1;
wire na673_1_i;
wire na674_1;
wire na674_1_i;
wire na675_1;
wire na675_1_i;
wire na676_1;
wire na676_1_i;
wire na677_1;
wire na677_1_i;
wire na678_1;
wire na678_1_i;
wire na679_1;
wire na679_1_i;
wire na680_1;
wire na680_1_i;
wire na681_1;
wire na681_1_i;
wire na682_1;
wire na682_1_i;
wire na683_1;
wire na683_1_i;
wire na684_1;
wire na684_1_i;
wire na685_1;
wire na685_1_i;
wire na686_1;
wire na686_1_i;
wire na687_1;
wire na687_1_i;
wire na688_1;
wire na688_1_i;
wire na689_1;
wire na689_1_i;
wire na690_1;
wire na690_1_i;
wire na691_1;
wire na691_1_i;
wire na692_1;
wire na692_1_i;
wire na693_1;
wire na693_1_i;
wire na694_1;
wire na694_1_i;
wire na695_1;
wire na695_1_i;
wire na696_1;
wire na696_1_i;
wire na697_1;
wire na697_1_i;
wire na698_1;
wire na698_1_i;
wire na699_1;
wire na699_1_i;
wire na700_1;
wire na700_1_i;
wire na701_1;
wire na701_1_i;
wire na702_1;
wire na702_1_i;
wire na703_1;
wire na703_1_i;
wire na704_1;
wire na704_1_i;
wire na705_1;
wire na705_1_i;
wire na706_1;
wire na706_1_i;
wire na707_1;
wire na707_1_i;
wire na708_1;
wire na708_1_i;
wire na709_1;
wire na709_1_i;
wire na710_1;
wire na710_1_i;
wire na711_1;
wire na711_1_i;
wire na712_1;
wire na712_1_i;
wire na713_1;
wire na713_1_i;
wire na714_1;
wire na714_1_i;
wire na715_1;
wire na715_1_i;
wire na716_1;
wire na716_1_i;
wire na717_1;
wire na717_1_i;
wire na718_1;
wire na718_1_i;
wire na719_1;
wire na719_1_i;
wire na720_1;
wire na720_1_i;
wire na721_1;
wire na721_1_i;
wire na722_1;
wire na722_1_i;
wire na723_1;
wire na723_1_i;
wire na724_1;
wire na724_1_i;
wire na725_1;
wire na725_1_i;
wire na726_1;
wire na726_1_i;
wire na727_1;
wire na727_1_i;
wire na728_1;
wire na728_1_i;
wire na729_1;
wire na729_1_i;
wire na730_1;
wire na730_1_i;
wire na731_1;
wire na731_1_i;
wire na732_1;
wire na732_1_i;
wire na733_1;
wire na733_1_i;
wire na734_1;
wire na734_1_i;
wire na735_1;
wire na735_1_i;
wire na736_1;
wire na736_1_i;
wire na737_1;
wire na737_1_i;
wire na738_1;
wire na738_1_i;
wire na739_1;
wire na739_1_i;
wire na740_1;
wire na740_1_i;
wire na741_1;
wire na741_1_i;
wire na742_1;
wire na742_1_i;
wire na743_1;
wire na743_1_i;
wire na744_1;
wire na744_1_i;
wire na745_1;
wire na745_1_i;
wire na746_1;
wire na746_1_i;
wire na747_1;
wire na747_1_i;
wire na748_1;
wire na748_1_i;
wire na749_1;
wire na749_1_i;
wire na750_1;
wire na750_1_i;
wire na751_1;
wire na751_1_i;
wire na752_1;
wire na752_1_i;
wire na753_1;
wire na753_1_i;
wire na754_1;
wire na754_1_i;
wire na755_1;
wire na755_1_i;
wire na756_1;
wire na756_1_i;
wire na757_1;
wire na757_1_i;
wire na758_1;
wire na758_1_i;
wire na759_1;
wire na759_1_i;
wire na760_1;
wire na760_1_i;
wire na761_1;
wire na761_1_i;
wire na762_1;
wire na762_1_i;
wire na763_1;
wire na763_1_i;
wire na764_1;
wire na764_1_i;
wire na765_1;
wire na765_1_i;
wire na766_1;
wire na766_1_i;
wire na767_1;
wire na767_1_i;
wire na768_1;
wire na768_1_i;
wire na769_1;
wire na769_1_i;
wire na770_1;
wire na770_1_i;
wire na771_1;
wire na771_1_i;
wire na772_1;
wire na772_1_i;
wire na773_1;
wire na773_1_i;
wire na774_1;
wire na774_1_i;
wire na775_1;
wire na775_1_i;
wire na776_1;
wire na776_1_i;
wire na777_1;
wire na777_1_i;
wire na778_1;
wire na778_1_i;
wire na779_1;
wire na779_1_i;
wire na780_1;
wire na780_1_i;
wire na781_1;
wire na781_1_i;
wire na782_1;
wire na782_1_i;
wire na783_1;
wire na783_1_i;
wire na784_1;
wire na784_1_i;
wire na785_1;
wire na785_1_i;
wire na786_1;
wire na786_1_i;
wire na787_1;
wire na787_1_i;
wire na788_1;
wire na788_1_i;
wire na789_1;
wire na789_1_i;
wire na790_1;
wire na790_1_i;
wire na791_1;
wire na791_1_i;
wire na792_1;
wire na792_1_i;
wire na793_1;
wire na793_1_i;
wire na794_1;
wire na794_1_i;
wire na795_1;
wire na795_1_i;
wire na796_1;
wire na796_1_i;
wire na797_1;
wire na797_1_i;
wire na798_1;
wire na798_1_i;
wire na799_1;
wire na799_1_i;
wire na800_1;
wire na800_1_i;
wire na801_1;
wire na801_1_i;
wire na802_1;
wire na802_1_i;
wire na803_1;
wire na803_1_i;
wire na804_1;
wire na804_1_i;
wire na805_1;
wire na805_1_i;
wire na806_1;
wire na806_1_i;
wire na807_1;
wire na807_1_i;
wire na808_2;
wire na808_2_i;
wire na809_1;
wire na809_2;
wire na810_2;
wire na810_2_i;
wire na811_1;
wire na811_1_i;
wire na812_1;
wire na812_1_i;
wire na813_1;
wire na813_1_i;
wire na814_2;
wire na814_2_i;
wire na815_1;
wire na815_1_i;
wire na816_1;
wire na816_2;
wire na817_1;
wire na818_2;
wire na819_1;
wire na820_1;
wire na821_1;
wire na821_2;
wire na822_2;
wire na824_1;
wire na824_2;
wire na825_1;
wire na826_1;
wire na827_1;
wire na827_2;
wire na829_1;
wire na832_1;
wire na834_1;
wire na836_1;
wire na838_1;
wire na839_1;
wire na842_2;
wire na843_1;
wire na844_1;
wire na845_1;
wire na846_2;
wire na848_1;
wire na849_1;
wire na850_1;
wire na851_1;
wire na852_1;
wire na853_1;
wire na854_1;
wire na855_2;
wire na857_1;
wire na858_1;
wire na859_1;
wire na860_1;
wire na861_1;
wire na861_1_i;
wire na862_1;
wire na862_2;
wire na863_2;
wire na864_2;
wire na865_1;
wire na866_1;
wire na867_2;
wire na868_1;
wire na869_1;
wire na870_1;
wire na870_1_i;
wire na871_1;
wire na871_2;
wire na872_1;
wire na873_2;
wire na874_1;
wire na875_1;
wire na876_1;
wire na876_1_i;
wire na877_1;
wire na877_2;
wire na878_1;
wire na880_1;
wire na881_1;
wire na882_1;
wire na882_1_i;
wire na883_1;
wire na883_2;
wire na884_2;
wire na886_1;
wire na886_1_i;
wire na887_1;
wire na887_2;
wire na888_1;
wire na889_1;
wire na889_1_i;
wire na890_1;
wire na890_2;
wire na891_1;
wire na891_1_i;
wire na892_1;
wire na892_2;
wire na893_2;
wire na894_1;
wire na894_1_i;
wire na895_1;
wire na895_2;
wire na896_1;
wire na897_1;
wire na898_1;
wire na899_2;
wire na900_1;
wire na901_1;
wire na901_2;
wire na903_1;
wire na903_2;
wire na904_1;
wire na906_1;
wire na909_1;
wire na911_1;
wire na913_1;
wire na914_1;
wire na915_2;
wire na916_1;
wire na917_1;
wire na919_1;
wire na920_1;
wire na921_1;
wire na925_1;
wire na926_1;
wire na927_1;
wire na929_1;
wire na929_2;
wire na930_1;
wire na932_1;
wire na933_2;
wire na934_1;
wire na935_1;
wire na936_1;
wire na937_1;
wire na938_1;
wire na939_1;
wire na939_1_i;
wire na940_1;
wire na940_2;
wire na942_1;
wire na943_1;
wire na944_1;
wire na945_1;
wire na946_1;
wire na947_1;
wire na948_1;
wire na948_1_i;
wire na949_1;
wire na949_2;
wire na950_1;
wire na951_1;
wire na952_1;
wire na953_2;
wire na954_1;
wire na954_1_i;
wire na955_1;
wire na955_2;
wire na956_1;
wire na957_2;
wire na958_2;
wire na959_1;
wire na960_1;
wire na961_1;
wire na961_1_i;
wire na962_1;
wire na962_2;
wire na963_1;
wire na964_1;
wire na964_1_i;
wire na965_1;
wire na965_2;
wire na966_2;
wire na967_1;
wire na967_1_i;
wire na968_1;
wire na968_2;
wire na969_1;
wire na969_1_i;
wire na970_1;
wire na970_2;
wire na971_1;
wire na971_1_i;
wire na972_1;
wire na972_2;
wire na973_1;
wire na975_2;
wire na976_1;
wire na977_1;
wire na977_2;
wire na978_2;
wire na979_1;
wire na979_2;
wire na981_1;
wire na981_2;
wire na982_1;
wire na984_1;
wire na987_2;
wire na989_1;
wire na991_1;
wire na992_1;
wire na993_1;
wire na994_1;
wire na995_1;
wire na996_1;
wire na997_1;
wire na998_1;
wire na999_1;
wire reset_n;
wire data_out;
wire na1000_1;
wire na1001_2;
wire na1002_2;
wire na1003_1;
wire na1004_1;
wire na1005_2;
wire na1006_1;
wire na1007_1;
wire na1008_1;
wire na1009_1;
wire na1010_1;
wire na1011_1;
wire na1012_1;
wire na1013_2;
wire na1014_1;
wire na1015_1;
wire na1016_1;
wire na1017_1;
wire na1017_1_i;
wire na1018_1;
wire na1018_2;
wire na1019_1;
wire na1022_2;
wire na1023_2;
wire na1024_1;
wire na1025_1;
wire na1026_1;
wire na1027_1;
wire na1028_1;
wire na1029_1;
wire na1029_1_i;
wire na1030_1;
wire na1030_2;
wire na1031_1;
wire na1032_1;
wire na1033_1;
wire na1034_1;
wire na1034_1_i;
wire na1035_1;
wire na1035_2;
wire na1036_1;
wire na1038_1;
wire na1039_1;
wire na1040_1;
wire na1040_1_i;
wire na1041_1;
wire na1041_2;
wire na1042_2;
wire na1044_1;
wire na1044_1_i;
wire na1045_1;
wire na1045_2;
wire na1046_1;
wire na1047_1;
wire na1048_1;
wire na1048_1_i;
wire na1049_1;
wire na1049_2;
wire na1050_1;
wire na1050_1_i;
wire na1051_1;
wire na1051_2;
wire na1052_1;
wire na1052_1_i;
wire na1053_1;
wire na1053_1_i;
wire na1054_1;
wire na1054_1_i;
wire na1055_1;
wire na1055_1_i;
wire na1056_1;
wire na1056_1_i;
wire na1057_1;
wire na1057_1_i;
wire na1058_1;
wire na1058_1_i;
wire na1059_1;
wire na1059_1_i;
wire na1060_1;
wire na1060_1_i;
wire na1061_1;
wire na1061_1_i;
wire na1062_1;
wire na1062_1_i;
wire na1063_1;
wire na1063_1_i;
wire na1064_1;
wire na1064_1_i;
wire na1065_1;
wire na1065_1_i;
wire na1066_1;
wire na1066_1_i;
wire na1067_1;
wire na1067_1_i;
wire na1068_1;
wire na1068_1_i;
wire na1069_1;
wire na1069_1_i;
wire na1070_1;
wire na1070_1_i;
wire na1071_1;
wire na1071_1_i;
wire na1072_1;
wire na1072_1_i;
wire na1073_1;
wire na1073_1_i;
wire na1074_1;
wire na1074_1_i;
wire na1075_1;
wire na1075_1_i;
wire na1076_1;
wire na1076_1_i;
wire na1077_1;
wire na1077_1_i;
wire na1078_1;
wire na1078_1_i;
wire na1079_1;
wire na1079_1_i;
wire na1080_1;
wire na1080_1_i;
wire na1081_1;
wire na1081_1_i;
wire na1082_1;
wire na1082_1_i;
wire na1083_1;
wire na1083_1_i;
wire na1084_1;
wire na1084_1_i;
wire na1085_1;
wire na1085_1_i;
wire na1086_1;
wire na1086_1_i;
wire na1087_1;
wire na1087_1_i;
wire na1088_1;
wire na1088_1_i;
wire na1089_1;
wire na1089_1_i;
wire na1090_1;
wire na1090_1_i;
wire na1091_1;
wire na1091_1_i;
wire na1092_1;
wire na1092_1_i;
wire na1093_1;
wire na1093_1_i;
wire na1094_1;
wire na1094_1_i;
wire na1095_1;
wire na1095_1_i;
wire na1096_1;
wire na1096_1_i;
wire na1097_1;
wire na1097_1_i;
wire na1098_1;
wire na1098_1_i;
wire na1099_1;
wire na1099_1_i;
wire na1100_1;
wire na1100_1_i;
wire na1101_1;
wire na1101_1_i;
wire na1102_1;
wire na1102_1_i;
wire na1103_1;
wire na1103_1_i;
wire na1104_1;
wire na1104_1_i;
wire na1105_1;
wire na1105_1_i;
wire na1106_1;
wire na1106_1_i;
wire na1107_1;
wire na1107_1_i;
wire na1108_1;
wire na1108_1_i;
wire na1109_1;
wire na1109_1_i;
wire na1110_1;
wire na1110_1_i;
wire na1111_1;
wire na1111_1_i;
wire na1112_1;
wire na1112_1_i;
wire na1113_1;
wire na1113_1_i;
wire na1114_1;
wire na1114_1_i;
wire na1115_1;
wire na1115_1_i;
wire na1116_1;
wire na1116_1_i;
wire na1117_1;
wire na1117_1_i;
wire na1118_1;
wire na1118_1_i;
wire na1119_1;
wire na1119_1_i;
wire na1120_1;
wire na1120_1_i;
wire na1121_1;
wire na1121_1_i;
wire na1122_1;
wire na1122_1_i;
wire na1123_1;
wire na1123_1_i;
wire na1124_1;
wire na1124_1_i;
wire na1125_1;
wire na1125_1_i;
wire na1126_1;
wire na1126_1_i;
wire na1127_1;
wire na1127_1_i;
wire na1128_1;
wire na1128_1_i;
wire na1129_1;
wire na1129_1_i;
wire na1130_1;
wire na1130_1_i;
wire na1131_1;
wire na1131_1_i;
wire na1132_1;
wire na1132_1_i;
wire na1133_1;
wire na1133_1_i;
wire na1134_1;
wire na1134_1_i;
wire na1135_1;
wire na1135_1_i;
wire na1136_1;
wire na1136_1_i;
wire na1137_1;
wire na1137_1_i;
wire na1138_1;
wire na1138_1_i;
wire na1139_1;
wire na1139_1_i;
wire na1140_1;
wire na1140_1_i;
wire na1141_1;
wire na1141_2;
wire na1142_1;
wire na1143_1;
wire na1143_2;
wire na1144_1;
wire na1144_2;
wire na1145_1;
wire na1145_2;
wire na1146_1;
wire na1146_2;
wire na1147_1;
wire na1147_2;
wire na1148_1;
wire na1148_2;
wire na1149_1;
wire na1149_2;
wire na1150_2;
wire na1150_2_i;
wire na1151_1;
wire na1151_1_i;
wire na1153_1;
wire na1154_1;
wire na1154_1_i;
wire na1155_1;
wire na1156_1;
wire na1156_1_i;
wire na1157_1;
wire na1158_1;
wire na1158_1_i;
wire na1159_1;
wire na1160_1;
wire na1160_1_i;
wire na1161_1;
wire na1162_1;
wire na1162_1_i;
wire na1163_1;
wire na1164_1;
wire na1164_1_i;
wire na1165_1;
wire na1166_1;
wire na1166_1_i;
wire na1167_1;
wire na1168_1;
wire na1168_1_i;
wire na1169_1;
wire na1170_1;
wire na1170_1_i;
wire na1171_1;
wire na1172_1;
wire na1172_1_i;
wire na1173_1;
wire na1174_1;
wire na1174_1_i;
wire na1175_1;
wire na1176_1;
wire na1176_1_i;
wire na1177_1;
wire na1178_1;
wire na1178_1_i;
wire na1179_1;
wire na1180_1;
wire na1180_1_i;
wire na1181_1;
wire na1182_1;
wire na1182_1_i;
wire na1183_1;
wire na1184_1;
wire na1184_1_i;
wire na1185_1;
wire na1186_1;
wire na1186_1_i;
wire na1187_1;
wire na1188_1;
wire na1188_1_i;
wire na1189_1;
wire na1190_1;
wire na1190_1_i;
wire na1191_1;
wire na1192_1;
wire na1192_1_i;
wire na1193_1;
wire na1194_1;
wire na1194_1_i;
wire na1195_1;
wire na1196_1;
wire na1196_1_i;
wire na1197_1;
wire na1198_1;
wire na1198_1_i;
wire na1199_1;
wire na1200_1;
wire na1200_1_i;
wire na1201_1;
wire na1202_1;
wire na1202_1_i;
wire na1203_1;
wire na1204_1;
wire na1204_1_i;
wire na1205_1;
wire na1206_1;
wire na1206_1_i;
wire na1207_1;
wire na1208_1;
wire na1208_1_i;
wire na1209_1;
wire na1210_1;
wire na1210_1_i;
wire na1211_1;
wire na1212_1;
wire na1212_1_i;
wire na1213_1;
wire na1214_1;
wire na1214_1_i;
wire na1215_1;
wire na1216_2;
wire na1216_2_i;
wire na1217_1;
wire na1217_1_i;
wire na1217_2;
wire na1217_2_i;
wire na1219_1;
wire na1219_1_i;
wire na1222_2;
wire na1223_1;
wire na1224_1;
wire na1224_2;
wire na1225_2;
wire na1228_1;
wire na1229_1;
wire na1230_1;
wire na1233_1;
wire na1235_1;
wire na1235_2;
wire na1236_1;
wire na1236_2;
wire na1238_2;
wire na1239_1;
wire na1243_1;
wire na1243_2;
wire na1245_1;
wire na1245_2;
wire na1246_2;
wire na1251_1;
wire na1251_2;
wire na1253_1;
wire na1253_1_i;
wire na1258_2;
wire na1259_1;
wire na1263_1;
wire na1265_1;
wire na1265_1_i;
wire na1270_1;
wire na1271_1;
wire na1277_1;
wire na1277_2;
wire na1280_1;
wire na1283_1;
wire na1286_1;
wire na1286_1_i;
wire na1289_1;
wire na1291_1;
wire na1291_2;
wire na1293_2;
wire na1294_1;
wire na1297_1;
wire na1297_1_i;
wire na1302_2;
wire na1303_1;
wire na1308_1;
wire na1308_1_i;
wire na1310_1;
wire na1313_1;
wire na1313_2;
wire na1315_1;
wire na1316_2;
wire na1319_1;
wire na1319_1_i;
wire na1323_1;
wire na1323_2;
wire na1325_1;
wire na1326_1;
wire na1331_1;
wire na1331_1_i;
wire na1332_1;
wire na1332_1_i;
wire na1333_1;
wire na1333_2;
wire na1335_1;
wire na1335_1_i;
wire na1335_2;
wire na1335_2_i;
wire na1336_2;
wire na1336_2_i;
wire na1337_1;
wire na1337_1_i;
wire na1338_2;
wire na1339_1;
wire na1342_1;
wire na1343_1;
wire na1343_1_i;
wire na1343_2;
wire na1343_2_i;
wire na1345_1;
wire na1345_1_i;
wire na1346_1;
wire na1346_1_i;
wire na1347_1;
wire na1348_1;
wire na1350_2;
wire na1351_1;
wire na1351_1_i;
wire na1353_2;
wire na1353_2_i;
wire na1355_1;
wire na1355_1_i;
wire na1355_2;
wire na1355_2_i;
wire na1356_2;
wire na1356_2_i;
wire na1357_2;
wire na1357_2_i;
wire na1358_1;
wire na1358_1_i;
wire na1358_2;
wire na1358_2_i;
wire na1359_1;
wire na1359_1_i;
wire na1359_2;
wire na1359_2_i;
wire na1361_1;
wire na1361_1_i;
wire na1362_1;
wire na1362_1_i;
wire na1363_1;
wire na1363_1_i;
wire na1364_1;
wire na1364_1_i;
wire na1365_1;
wire na1365_1_i;
wire na1366_1;
wire na1366_1_i;
wire na1367_1;
wire na1367_1_i;
wire na1368_1;
wire na1368_1_i;
wire na1369_1;
wire na1369_1_i;
wire na1370_2;
wire na1370_2_i;
wire na1371_1;
wire na1372_1;
wire na1375_1;
wire na1376_1;
wire na1376_1_i;
wire na1377_1;
wire na1377_1_i;
wire na1377_2;
wire na1377_2_i;
wire na1378_1;
wire na1378_1_i;
wire na1379_1;
wire na1379_1_i;
wire na1379_2;
wire na1379_2_i;
wire na1380_1;
wire na1380_1_i;
wire na1382_2;
wire na1382_2_i;
wire na1383_1;
wire na1383_1_i;
wire na1383_2;
wire na1383_2_i;
wire na1386_2;
wire na1386_2_i;
wire na1387_1;
wire na1387_2;
wire na1388_2;
wire na1389_1;
wire na1390_2;
wire na1391_1;
wire na1392_2;
wire na1393_1;
wire na1394_1;
wire na1395_1;
wire na1396_1;
wire na1397_2;
wire na1398_1;
wire na1399_2;
wire na1400_1;
wire na1401_2;
wire na1402_1;
wire na1403_2;
wire na1404_1;
wire na1405_1;
wire na1406_2;
wire na1407_2;
wire na1408_1;
wire na1409_1;
wire na1410_2;
wire na1411_1;
wire na1412_1;
wire na1413_2;
wire na1414_2;
wire na1415_2;
wire na1416_2;
wire na1417_1;
wire na1418_1;
wire na1419_1;
wire na1420_1;
wire na1421_2;
wire na1422_1;
wire na1423_1;
wire na1424_1;
wire na1425_2;
wire na1426_2;
wire na1427_1;
wire na1428_2;
wire na1429_1;
wire na1430_2;
wire na1431_2;
wire na1432_1;
wire na1433_1;
wire na1434_2;
wire na1435_2;
wire na1436_1;
wire na1437_2;
wire na1438_2;
wire na1439_1;
wire na1440_2;
wire na1441_2;
wire na1442_1;
wire na1443_1;
wire na1444_1;
wire na1445_2;
wire na1446_1;
wire na1447_1;
wire na1448_2;
wire na1449_1;
wire na1450_2;
wire na1451_1;
wire na1451_2;
wire na1452_1;
wire na1453_1;
wire na1454_1;
wire na1455_1;
wire na1456_2;
wire na1458_1;
wire na1459_1;
wire na1460_2;
wire na1461_1;
wire na1462_1;
wire na1463_2;
wire na1464_1;
wire na1465_1;
wire na1466_1;
wire na1467_2;
wire na1468_1;
wire na1469_1;
wire na1470_2;
wire na1471_2;
wire na1472_1;
wire na1473_1;
wire na1474_1;
wire na1475_1;
wire na1477_2;
wire na1478_1;
wire na1479_2;
wire na1480_2;
wire na1481_1;
wire na1482_1;
wire na1482_2;
wire na1483_1;
wire na1483_2;
wire na1484_1;
wire na1484_2;
wire na1486_1;
wire na1486_2;
wire na1488_1;
wire na1488_2;
wire na1490_1;
wire na1490_2;
wire na1492_1;
wire na1492_2;
wire na1493_1;
wire na1493_2;
wire na1494_1;
wire na1494_2;
wire na1495_2;
wire na1495_2_i;
wire na1496_1;
wire na1496_1_i;
wire na1497_1;
wire na1497_1_i;
wire na1498_1;
wire na1498_1_i;
wire na1499_1;
wire na1499_2;
wire na1500_1;
wire na1500_2;
wire na1501_2;
wire na1501_2_i;
wire na1502_1;
wire na1502_2;
wire na1503_1;
wire na1503_1_i;
wire na1504_1;
wire na1504_2;
wire na1505_2;
wire na1505_2_i;
wire na1506_2;
wire na1506_2_i;
wire na1507_1;
wire na1507_2;
wire na1508_1;
wire na1508_2;
wire na1509_1;
wire na1509_2;
wire na1510_2;
wire na1510_2_i;
wire na1511_1;
wire na1511_1_i;
wire na1512_1;
wire na1512_2;
wire na1513_1;
wire na1513_2;
wire na1514_1;
wire na1514_1_i;
wire na1515_1;
wire na1515_1_i;
wire na1516_1;
wire na1516_2;
wire na1517_2;
wire na1517_2_i;
wire na1518_2;
wire na1518_2_i;
wire na1519_2;
wire na1519_2_i;
wire na1520_1;
wire na1520_1_i;
wire na1521_2;
wire na1521_2_i;
wire na1522_2;
wire na1522_2_i;
wire na1523_2;
wire na1523_2_i;
wire na1524_1;
wire na1524_1_i;
wire na1525_2;
wire na1525_2_i;
wire na1526_1;
wire na1526_1_i;
wire na1527_1;
wire na1527_1_i;
wire na1528_1;
wire na1528_1_i;
wire na1529_1;
wire na1529_2;
wire na1530_1;
wire na1530_2;
wire na1531_2;
wire na1531_2_i;
wire na1532_2;
wire na1532_2_i;
wire na1533_2;
wire na1533_2_i;
wire na1534_2;
wire na1534_2_i;
wire na1535_2;
wire na1535_2_i;
wire na1536_1;
wire na1536_1_i;
wire na1537_1;
wire na1537_1_i;
wire na1538_1;
wire na1538_2;
wire na1539_1;
wire na1539_2;
wire na1540_1;
wire na1540_1_i;
wire na1541_1;
wire na1541_2;
wire na1542_2;
wire na1542_2_i;
wire na1543_2;
wire na1543_2_i;
wire na1544_2;
wire na1544_2_i;
wire na1545_1;
wire na1545_1_i;
wire na1546_2;
wire na1546_2_i;
wire na1547_1;
wire na1547_1_i;
wire na1548_1;
wire na1548_1_i;
wire na1549_1;
wire na1549_1_i;
wire na1550_1;
wire na1550_1_i;
wire na1551_1;
wire na1551_1_i;
wire na1552_2;
wire na1552_2_i;
wire na1553_1;
wire na1553_1_i;
wire na1554_1;
wire na1554_1_i;
wire na1555_2;
wire na1555_2_i;
wire na1556_1;
wire na1556_1_i;
wire na1557_1;
wire na1557_1_i;
wire na1558_2;
wire na1558_2_i;
wire na1559_1;
wire na1559_1_i;
wire na1560_1;
wire na1560_1_i;
wire na1561_2;
wire na1561_2_i;
wire na1562_2;
wire na1562_2_i;
wire na1563_2;
wire na1563_2_i;
wire na1564_1;
wire na1564_1_i;
wire na1565_2;
wire na1565_2_i;
wire na1566_2;
wire na1566_2_i;
wire na1567_1;
wire na1567_1_i;
wire na1568_1;
wire na1568_1_i;
wire na1569_2;
wire na1569_2_i;
wire na1570_2;
wire na1570_2_i;
wire na1571_1;
wire na1571_1_i;
wire na1572_2;
wire na1572_2_i;
wire na1573_1;
wire na1573_1_i;
wire na1574_1;
wire na1574_1_i;
wire na1575_2;
wire na1575_2_i;
wire na1576_1;
wire na1576_1_i;
wire na1577_2;
wire na1577_2_i;
wire na1578_1;
wire na1578_1_i;
wire na1579_2;
wire na1579_2_i;
wire na1580_1;
wire na1580_1_i;
wire na1581_2;
wire na1581_2_i;
wire na1582_2;
wire na1582_2_i;
wire na1583_1;
wire na1583_1_i;
wire na1584_1;
wire na1584_1_i;
wire na1585_1;
wire na1585_1_i;
wire na1586_1;
wire na1586_1_i;
wire na1587_2;
wire na1587_2_i;
wire na1588_2;
wire na1588_2_i;
wire na1589_1;
wire na1589_1_i;
wire na1590_2;
wire na1590_2_i;
wire na1591_1;
wire na1591_1_i;
wire na1592_1;
wire na1592_1_i;
wire na1593_1;
wire na1593_1_i;
wire na1594_1;
wire na1594_1_i;
wire na1595_2;
wire na1595_2_i;
wire na1596_1;
wire na1596_1_i;
wire na1597_2;
wire na1597_2_i;
wire na1598_1;
wire na1598_1_i;
wire na1599_1;
wire na1599_1_i;
wire na1600_1;
wire na1600_1_i;
wire na1601_2;
wire na1601_2_i;
wire na1602_2;
wire na1602_2_i;
wire na1603_2;
wire na1603_2_i;
wire na1604_2;
wire na1604_2_i;
wire na1605_1;
wire na1605_1_i;
wire na1606_2;
wire na1606_2_i;
wire na1607_1;
wire na1607_1_i;
wire na1608_2;
wire na1608_2_i;
wire na1609_1;
wire na1609_1_i;
wire na1610_2;
wire na1610_2_i;
wire na1611_2;
wire na1611_2_i;
wire na1612_1;
wire na1612_1_i;
wire na1613_2;
wire na1613_2_i;
wire na1614_1;
wire na1614_2;
wire na1615_1;
wire na1615_1_i;
wire na1616_2;
wire na1616_2_i;
wire na1617_1;
wire na1617_1_i;
wire na1618_2;
wire na1618_2_i;
wire na1619_1;
wire na1619_2;
wire na1620_1;
wire na1620_2;
wire na1621_2;
wire na1621_2_i;
wire na1622_1;
wire na1622_2;
wire na1623_2;
wire na1623_2_i;
wire na1624_1;
wire na1624_2;
wire na1625_1;
wire na1625_1_i;
wire na1626_1;
wire na1626_1_i;
wire na1627_1;
wire na1627_2;
wire na1628_1;
wire na1628_2;
wire na1629_1;
wire na1629_2;
wire na1630_1;
wire na1630_1_i;
wire na1631_2;
wire na1631_2_i;
wire na1632_1;
wire na1632_2;
wire na1633_1;
wire na1633_2;
wire na1634_2;
wire na1634_2_i;
wire na1635_2;
wire na1635_2_i;
wire na1636_1;
wire na1636_2;
wire na1637_1;
wire na1637_1_i;
wire na1638_1;
wire na1638_2;
wire na1639_1;
wire na1639_2;
wire na1640_1;
wire na1640_2;
wire na1641_1;
wire na1641_2;
wire na1642_1;
wire na1642_2;
wire na1643_1;
wire na1643_2;
wire na1644_2;
wire na1644_2_i;
wire na1645_1;
wire na1645_1_i;
wire na1646_1;
wire na1646_1_i;
wire na1647_2;
wire na1647_2_i;
wire na1648_1;
wire na1648_1_i;
wire na1649_2;
wire na1649_2_i;
wire na1650_1;
wire na1650_1_i;
wire na1651_1;
wire na1651_1_i;
wire na1652_2;
wire na1652_2_i;
wire na1653_2;
wire na1653_2_i;
wire na1654_2;
wire na1654_2_i;
wire na1655_1;
wire na1655_1_i;
wire na1656_2;
wire na1656_2_i;
wire na1657_1;
wire na1657_2;
wire na1658_1;
wire na1658_2;
wire na1659_1;
wire na1659_1_i;
wire na1660_1;
wire na1660_1_i;
wire na1661_1;
wire na1661_1_i;
wire na1662_1;
wire na1662_1_i;
wire na1663_2;
wire na1663_2_i;
wire na1664_2;
wire na1664_2_i;
wire na1665_1;
wire na1665_1_i;
wire na1666_1;
wire na1666_2;
wire na1667_1;
wire na1667_2;
wire na1668_1;
wire na1668_1_i;
wire na1669_1;
wire na1669_2;
wire na1670_2;
wire na1670_2_i;
wire na1671_2;
wire na1671_2_i;
wire na1672_2;
wire na1672_2_i;
wire na1673_1;
wire na1673_1_i;
wire na1674_2;
wire na1674_2_i;
wire na1675_1;
wire na1675_1_i;
wire na1676_1;
wire na1676_2;
wire na1677_1;
wire na1677_2;
wire na1678_1;
wire na1678_1_i;
wire na1679_1;
wire na1679_1_i;
wire na1680_2;
wire na1680_2_i;
wire na1681_1;
wire na1681_1_i;
wire na1682_2;
wire na1682_2_i;
wire na1683_2;
wire na1683_2_i;
wire na1684_1;
wire na1684_1_i;
wire na1685_2;
wire na1685_2_i;
wire na1686_2;
wire na1686_2_i;
wire na1687_1;
wire na1687_1_i;
wire na1688_1;
wire na1688_1_i;
wire na1689_2;
wire na1689_2_i;
wire na1690_1;
wire na1690_1_i;
wire na1691_2;
wire na1691_2_i;
wire na1692_1;
wire na1692_1_i;
wire na1693_2;
wire na1693_2_i;
wire na1694_1;
wire na1694_1_i;
wire na1695_2;
wire na1695_2_i;
wire na1696_1;
wire na1696_1_i;
wire na1697_1;
wire na1697_1_i;
wire na1698_2;
wire na1698_2_i;
wire na1699_1;
wire na1699_1_i;
wire na1700_1;
wire na1700_1_i;
wire na1701_2;
wire na1701_2_i;
wire na1702_1;
wire na1702_1_i;
wire na1703_1;
wire na1703_1_i;
wire na1704_1;
wire na1704_1_i;
wire na1705_2;
wire na1705_2_i;
wire na1706_1;
wire na1706_1_i;
wire na1707_2;
wire na1707_2_i;
wire na1708_1;
wire na1708_1_i;
wire na1709_2;
wire na1709_2_i;
wire na1710_2;
wire na1710_2_i;
wire na1711_1;
wire na1711_1_i;
wire na1712_1;
wire na1712_1_i;
wire na1713_1;
wire na1713_1_i;
wire na1714_1;
wire na1714_1_i;
wire na1715_1;
wire na1715_1_i;
wire na1716_1;
wire na1716_1_i;
wire na1717_1;
wire na1717_1_i;
wire na1718_2;
wire na1718_2_i;
wire na1719_1;
wire na1719_1_i;
wire na1720_1;
wire na1720_1_i;
wire na1721_1;
wire na1721_1_i;
wire na1722_2;
wire na1722_2_i;
wire na1723_2;
wire na1723_2_i;
wire na1724_2;
wire na1724_2_i;
wire na1725_1;
wire na1725_1_i;
wire na1726_1;
wire na1726_1_i;
wire na1727_1;
wire na1727_1_i;
wire na1728_2;
wire na1728_2_i;
wire na1729_2;
wire na1729_2_i;
wire na1730_1;
wire na1730_1_i;
wire na1731_1;
wire na1731_1_i;
wire na1732_1;
wire na1732_1_i;
wire na1733_2;
wire na1733_2_i;
wire na1734_1;
wire na1734_1_i;
wire na1735_1;
wire na1735_1_i;
wire na1736_1;
wire na1736_1_i;
wire na1737_2;
wire na1737_2_i;
wire na1738_1;
wire na1738_1_i;
wire na1739_1;
wire na1739_1_i;
wire na1740_2;
wire na1740_2_i;
wire na1741_2;
wire na1741_2_i;
wire na1742_1;
wire na1743_2;
wire na1744_2;
wire na1745_2;
wire na1746_1;
wire na1747_1;
wire na1749_1;
wire na1751_1;
wire na1753_1;
wire na1755_1;
wire na1757_1;
wire na1759_1;
wire na1760_2;
wire na1761_2;
wire na1762_1;
wire na1764_1;
wire na1766_1;
wire na1768_1;
wire na1770_1;
wire na1772_1;
wire na1774_1;
wire na1775_1;
wire na1777_1;
wire na1779_1;
wire na1781_1;
wire na1783_1;
wire na1784_1;
wire na1785_1;
wire na1787_1;
wire na1789_1;
wire na1790_2;
wire na1791_1;
wire na1793_1;
wire na1795_1;
wire na1797_1;
wire na1798_1;
wire na1810_1;
wire na1811_1;
wire na1812_1;
wire na1813_1;
wire na1814_1;
wire na1816_1;
wire na1817_1;
wire na1818_1;
wire na1819_1;
wire na1819_1_i;
wire na1821_1;
wire na1822_2;
wire na1823_1;
wire na1824_1;
wire na1824_1_i;
wire na1826_1;
wire na1827_1;
wire na1828_1;
wire na1829_1;
wire na1829_1_i;
wire na1831_1;
wire na1832_1;
wire na1833_1;
wire na1834_1;
wire na1834_1_i;
wire na1835_2;
wire na1836_1;
wire na1837_1;
wire na1838_1;
wire na1838_1_i;
wire na1839_1;
wire na1840_2;
wire na1841_2;
wire na1842_1;
wire na1844_1;
wire na1845_1;
wire na1846_2;
wire na1847_2;
wire na1848_1;
wire na1850_1;
wire na1851_2;
wire na1852_1;
wire na1853_1;
wire na1855_1;
wire na1856_1;
wire na1857_1;
wire na1857_1_i;
wire na1858_1;
wire na1859_1;
wire na1859_1_i;
wire na1861_1;
wire na1862_1;
wire na1862_1_i;
wire na1864_4;
wire na1866_4;
wire na1868_4;
wire na1870_4;
wire na1871_1;
wire na1871_4;
wire na1872_1;
wire na1872_2;
wire na1872_4;
wire na1874_1;
wire na1874_2;
wire na1874_4;
wire na1876_1;
wire na1877_1;
wire na1877_4;
wire na1878_1;
wire na1878_2;
wire na1878_4;
wire na1880_1;
wire na1880_2;
wire na1882_1;
wire na1882_4;
wire na1883_1;
wire na1883_2;
wire na1883_4;
wire na1885_1;
wire na1886_1;
wire na1886_4;
wire na1888_1;
wire na1888_2;
wire na1888_4;
wire na1890_1;
wire na1890_2;
wire na1890_4;
wire na1892_1;
wire na1892_2;
wire na1892_4;
wire na1894_1;
wire na1894_2;
wire na1894_4;
wire na1896_1;
wire na1896_2;
wire na1897_1;
wire na1897_4;
wire na1898_1;
wire na1898_2;
wire na1900_1;
wire na1900_4;
wire na1902_1;
wire na1902_2;
wire na1902_4;
wire na1904_1;
wire na1904_2;
wire na1904_4;
wire na1906_1;
wire na1906_2;
wire na1906_4;
wire na1908_1;
wire na1908_2;
wire na1908_4;
wire na1910_1;
wire na1910_2;
wire na1911_1;
wire na1911_4;
wire na1912_1;
wire na1912_2;
wire na1915_1;
wire na1915_1_i;
wire na1916_2;
wire na1916_2_i;
wire na1917_1;
wire na1917_1_i;
wire na1918_2;
wire na1918_2_i;
wire na1919_1;
wire na1919_1_i;
wire na1920_2;
wire na1920_2_i;
wire na1921_2;
wire na1921_2_i;
wire na1922_1;
wire na1922_1_i;
wire na1923_1;
wire na1924_2;
wire na1924_2_i;
wire na1925_1;
wire na1925_1_i;
wire na1926_2;
wire na1926_2_i;
wire na1927_1;
wire na1927_1_i;
wire na1928_2;
wire na1928_2_i;
wire na1929_1;
wire na1929_1_i;
wire na1930_2;
wire na1930_2_i;
wire na1931_1;
wire na1931_1_i;
wire na1961_2;
wire na1961_2_i;
wire na1962_1;
wire na1962_1_i;
wire na1963_2;
wire na1963_2_i;
wire na1964_1;
wire na1964_1_i;
wire na1965_2;
wire na1965_2_i;
wire na1966_1;
wire na1966_1_i;
wire na1967_2;
wire na1967_2_i;
wire na1968_1;
wire na1968_1_i;
wire na1971_2;
wire na1971_2_i;
wire na1972_1;
wire na1972_1_i;
wire na1973_2;
wire na1973_2_i;
wire na1974_1;
wire na1974_1_i;
wire na1975_2;
wire na1975_2_i;
wire na1976_1;
wire na1976_1_i;
wire na1977_2;
wire na1977_2_i;
wire na1978_1;
wire na1978_1_i;
wire na1979_2;
wire na1979_2_i;
wire na1980_1;
wire na1980_1_i;
wire na1981_2;
wire na1981_2_i;
wire na1982_1;
wire na1982_1_i;
wire na1983_2;
wire na1983_2_i;
wire na1984_2;
wire na1984_2_i;
wire na1985_2;
wire na1985_2_i;
wire na1986_1;
wire na1986_1_i;
wire na1987_2;
wire na1987_2_i;
wire na1988_1;
wire na1988_1_i;
wire na1989_2;
wire na1989_2_i;
wire na1990_1;
wire na1990_1_i;
wire na1991_2;
wire na1991_2_i;
wire na1992_1;
wire na1992_1_i;
wire na1993_2;
wire na1993_2_i;
wire na1994_1;
wire na1994_1_i;
wire na1995_2;
wire na1995_2_i;
wire na1996_1;
wire na1996_1_i;
wire na1997_2;
wire na1997_2_i;
wire na1998_1;
wire na1998_1_i;
wire na1999_2;
wire na1999_2_i;
wire na2000_1;
wire na2000_1_i;
wire na2001_2;
wire na2001_2_i;
wire na2002_1;
wire na2002_1_i;
wire na2003_2;
wire na2003_2_i;
wire na2004_1;
wire na2004_1_i;
wire na2005_2;
wire na2005_2_i;
wire na2006_1;
wire na2006_1_i;
wire na2007_2;
wire na2007_2_i;
wire na2008_1;
wire na2008_1_i;
wire na2009_2;
wire na2009_2_i;
wire na2010_1;
wire na2010_1_i;
wire na2011_2;
wire na2011_2_i;
wire na2012_1;
wire na2012_1_i;
wire na2013_2;
wire na2013_2_i;
wire na2014_1;
wire na2014_1_i;
wire na2015_2;
wire na2015_2_i;
wire na2016_1;
wire na2016_1_i;
wire na2017_2;
wire na2017_2_i;
wire na2018_1;
wire na2018_1_i;
wire na2019_2;
wire na2019_2_i;
wire na2020_1;
wire na2020_1_i;
wire na2021_2;
wire na2021_2_i;
wire na2022_1;
wire na2022_1_i;
wire na2023_2;
wire na2023_2_i;
wire na2024_1;
wire na2024_1_i;
wire na2025_2;
wire na2025_2_i;
wire na2026_1;
wire na2026_1_i;
wire na2027_2;
wire na2027_2_i;
wire na2028_1;
wire na2028_1_i;
wire na2029_2;
wire na2029_2_i;
wire na2030_1;
wire na2030_1_i;
wire na2031_2;
wire na2031_2_i;
wire na2032_1;
wire na2032_1_i;
wire na2033_2;
wire na2033_2_i;
wire na2034_1;
wire na2034_1_i;
wire na2035_2;
wire na2035_2_i;
wire na2036_1;
wire na2036_1_i;
wire na2037_2;
wire na2037_2_i;
wire na2038_1;
wire na2038_1_i;
wire na2039_2;
wire na2039_2_i;
wire na2040_1;
wire na2040_1_i;
wire na2041_2;
wire na2041_2_i;
wire na2042_1;
wire na2042_1_i;
wire na2043_2;
wire na2043_2_i;
wire na2044_1;
wire na2044_1_i;
wire na2045_1;
wire na2045_1_i;
wire na2046_1;
wire na2046_1_i;
wire na2047_2;
wire na2047_2_i;
wire na2048_1;
wire na2048_1_i;
wire na2049_2;
wire na2049_2_i;
wire na2050_1;
wire na2050_1_i;
wire na2051_2;
wire na2051_2_i;
wire na2052_1;
wire na2052_1_i;
wire na2053_2;
wire na2053_2_i;
wire na2054_1;
wire na2054_1_i;
wire na2055_2;
wire na2055_2_i;
wire na2056_1;
wire na2056_1_i;
wire na2057_2;
wire na2057_2_i;
wire na2058_1;
wire na2058_1_i;
wire na2059_2;
wire na2059_2_i;
wire na2060_1;
wire na2060_1_i;
wire na2061_2;
wire na2061_2_i;
wire na2062_1;
wire na2062_1_i;
wire na2063_2;
wire na2063_2_i;
wire na2064_1;
wire na2064_1_i;
wire na2065_2;
wire na2065_2_i;
wire na2066_1;
wire na2066_1_i;
wire na2067_2;
wire na2067_2_i;
wire na2068_1;
wire na2068_1_i;
wire na2069_2;
wire na2069_2_i;
wire na2070_1;
wire na2070_1_i;
wire na2071_2;
wire na2071_2_i;
wire na2072_1;
wire na2072_1_i;
wire na2073_2;
wire na2073_2_i;
wire na2074_1;
wire na2074_1_i;
wire na2075_2;
wire na2075_2_i;
wire na2076_1;
wire na2076_1_i;
wire na2077_2;
wire na2077_2_i;
wire na2078_1;
wire na2078_1_i;
wire na2079_2;
wire na2079_2_i;
wire na2080_1;
wire na2080_1_i;
wire na2081_2;
wire na2081_2_i;
wire na2082_1;
wire na2082_1_i;
wire na2083_2;
wire na2083_2_i;
wire na2084_1;
wire na2084_1_i;
wire na2085_2;
wire na2085_2_i;
wire na2086_1;
wire na2086_1_i;
wire na2087_2;
wire na2087_2_i;
wire na2088_1;
wire na2088_1_i;
wire na2089_2;
wire na2089_2_i;
wire na2090_1;
wire na2090_1_i;
wire na2091_2;
wire na2091_2_i;
wire na2092_1;
wire na2092_1_i;
wire na2093_2;
wire na2093_2_i;
wire na2094_1;
wire na2094_1_i;
wire na2095_2;
wire na2095_2_i;
wire na2096_1;
wire na2096_1_i;
wire na2097_2;
wire na2097_2_i;
wire na2098_1;
wire na2098_1_i;
wire na2099_2;
wire na2099_2_i;
wire na2100_1;
wire na2100_1_i;
wire na2101_2;
wire na2101_2_i;
wire na2102_1;
wire na2102_1_i;
wire na2103_2;
wire na2103_2_i;
wire na2104_1;
wire na2104_1_i;
wire na2105_2;
wire na2105_2_i;
wire na2106_2;
wire na2106_2_i;
wire na2107_2;
wire na2107_2_i;
wire na2108_1;
wire na2108_1_i;
wire na2109_2;
wire na2109_2_i;
wire na2110_1;
wire na2110_1_i;
wire na2111_2;
wire na2111_2_i;
wire na2112_1;
wire na2112_1_i;
wire na2113_2;
wire na2113_2_i;
wire na2114_1;
wire na2114_1_i;
wire na2115_2;
wire na2115_2_i;
wire na2116_1;
wire na2116_1_i;
wire na2117_2;
wire na2117_2_i;
wire na2118_1;
wire na2118_1_i;
wire na2119_2;
wire na2119_2_i;
wire na2120_1;
wire na2120_1_i;
wire na2121_2;
wire na2121_2_i;
wire na2122_1;
wire na2122_1_i;
wire na2123_2;
wire na2123_2_i;
wire na2124_1;
wire na2124_1_i;
wire na2125_2;
wire na2125_2_i;
wire na2126_1;
wire na2126_1_i;
wire na2127_2;
wire na2127_2_i;
wire na2128_1;
wire na2128_1_i;
wire na2129_2;
wire na2129_2_i;
wire na2130_1;
wire na2130_1_i;
wire na2131_2;
wire na2131_2_i;
wire na2132_1;
wire na2132_1_i;
wire na2133_2;
wire na2133_2_i;
wire na2134_1;
wire na2134_1_i;
wire na2135_2;
wire na2135_2_i;
wire na2136_1;
wire na2136_1_i;
wire na2137_2;
wire na2137_2_i;
wire na2138_1;
wire na2138_1_i;
wire na2139_2;
wire na2139_2_i;
wire na2140_1;
wire na2140_1_i;
wire na2141_2;
wire na2141_2_i;
wire na2142_1;
wire na2142_1_i;
wire na2143_2;
wire na2143_2_i;
wire na2144_1;
wire na2144_1_i;
wire na2145_2;
wire na2145_2_i;
wire na2146_1;
wire na2146_1_i;
wire na2147_2;
wire na2147_2_i;
wire na2148_1;
wire na2148_1_i;
wire na2149_2;
wire na2149_2_i;
wire na2150_1;
wire na2150_1_i;
wire na2151_2;
wire na2151_2_i;
wire na2152_1;
wire na2152_1_i;
wire na2153_2;
wire na2153_2_i;
wire na2154_1;
wire na2154_1_i;
wire na2155_2;
wire na2155_2_i;
wire na2156_1;
wire na2156_1_i;
wire na2157_2;
wire na2157_2_i;
wire na2158_1;
wire na2158_1_i;
wire na2159_2;
wire na2159_2_i;
wire na2160_1;
wire na2160_1_i;
wire na2161_2;
wire na2161_2_i;
wire na2162_1;
wire na2162_1_i;
wire na2163_2;
wire na2163_2_i;
wire na2164_1;
wire na2164_1_i;
wire na2165_2;
wire na2165_2_i;
wire na2166_1;
wire na2166_1_i;
wire na2167_1;
wire na2167_1_i;
wire na2168_1;
wire na2168_1_i;
wire na2169_2;
wire na2169_2_i;
wire na2170_1;
wire na2170_1_i;
wire na2171_2;
wire na2171_2_i;
wire na2172_1;
wire na2172_1_i;
wire na2173_2;
wire na2173_2_i;
wire na2174_1;
wire na2174_1_i;
wire na2175_2;
wire na2175_2_i;
wire na2176_1;
wire na2176_1_i;
wire na2177_2;
wire na2177_2_i;
wire na2178_1;
wire na2178_1_i;
wire na2179_2;
wire na2179_2_i;
wire na2180_1;
wire na2180_1_i;
wire na2181_2;
wire na2181_2_i;
wire na2182_1;
wire na2182_1_i;
wire na2183_2;
wire na2183_2_i;
wire na2184_1;
wire na2184_1_i;
wire na2185_2;
wire na2185_2_i;
wire na2186_1;
wire na2186_1_i;
wire na2187_2;
wire na2187_2_i;
wire na2188_1;
wire na2188_1_i;
wire na2189_2;
wire na2189_2_i;
wire na2190_1;
wire na2190_1_i;
wire na2191_2;
wire na2191_2_i;
wire na2192_1;
wire na2192_1_i;
wire na2193_2;
wire na2193_2_i;
wire na2194_1;
wire na2194_1_i;
wire na2195_2;
wire na2195_2_i;
wire na2196_1;
wire na2196_1_i;
wire na2197_2;
wire na2197_2_i;
wire na2198_1;
wire na2198_1_i;
wire na2199_2;
wire na2199_2_i;
wire na2200_1;
wire na2200_1_i;
wire na2201_2;
wire na2201_2_i;
wire na2202_1;
wire na2202_1_i;
wire na2203_2;
wire na2203_2_i;
wire na2204_1;
wire na2204_1_i;
wire na2205_2;
wire na2205_2_i;
wire na2206_1;
wire na2206_1_i;
wire na2207_2;
wire na2207_2_i;
wire na2208_1;
wire na2208_1_i;
wire na2209_2;
wire na2209_2_i;
wire na2210_1;
wire na2210_1_i;
wire na2211_2;
wire na2211_2_i;
wire na2212_1;
wire na2212_1_i;
wire na2213_2;
wire na2213_2_i;
wire na2214_1;
wire na2214_1_i;
wire na2215_2;
wire na2215_2_i;
wire na2216_1;
wire na2216_1_i;
wire na2217_2;
wire na2217_2_i;
wire na2218_1;
wire na2218_1_i;
wire na2219_2;
wire na2219_2_i;
wire na2220_1;
wire na2220_1_i;
wire na2221_2;
wire na2221_2_i;
wire na2222_1;
wire na2222_1_i;
wire na2223_2;
wire na2223_2_i;
wire na2224_1;
wire na2224_1_i;
wire na2225_2;
wire na2225_2_i;
wire na2226_1;
wire na2226_1_i;
wire na2227_2;
wire na2227_2_i;
wire na2228_2;
wire na2228_2_i;
wire na2229_2;
wire na2229_2_i;
wire na2230_1;
wire na2230_1_i;
wire na2231_2;
wire na2231_2_i;
wire na2232_1;
wire na2232_1_i;
wire na2233_2;
wire na2233_2_i;
wire na2234_1;
wire na2234_1_i;
wire na2235_2;
wire na2235_2_i;
wire na2236_1;
wire na2236_1_i;
wire na2237_2;
wire na2237_2_i;
wire na2238_1;
wire na2238_1_i;
wire na2239_2;
wire na2239_2_i;
wire na2240_1;
wire na2240_1_i;
wire na2241_2;
wire na2241_2_i;
wire na2242_1;
wire na2242_1_i;
wire na2243_2;
wire na2243_2_i;
wire na2244_1;
wire na2244_1_i;
wire na2245_2;
wire na2245_2_i;
wire na2246_1;
wire na2246_1_i;
wire na2247_2;
wire na2247_2_i;
wire na2248_1;
wire na2248_1_i;
wire na2249_2;
wire na2249_2_i;
wire na2250_1;
wire na2250_1_i;
wire na2251_2;
wire na2251_2_i;
wire na2252_1;
wire na2252_1_i;
wire na2253_2;
wire na2253_2_i;
wire na2254_1;
wire na2254_1_i;
wire na2255_2;
wire na2255_2_i;
wire na2256_1;
wire na2256_1_i;
wire na2257_2;
wire na2257_2_i;
wire na2258_1;
wire na2258_1_i;
wire na2259_2;
wire na2259_2_i;
wire na2260_1;
wire na2260_1_i;
wire na2261_2;
wire na2261_2_i;
wire na2262_1;
wire na2262_1_i;
wire na2263_2;
wire na2263_2_i;
wire na2264_1;
wire na2264_1_i;
wire na2265_2;
wire na2265_2_i;
wire na2266_1;
wire na2266_1_i;
wire na2267_2;
wire na2267_2_i;
wire na2268_1;
wire na2268_1_i;
wire na2269_2;
wire na2269_2_i;
wire na2270_1;
wire na2270_1_i;
wire na2271_2;
wire na2271_2_i;
wire na2272_1;
wire na2272_1_i;
wire na2273_2;
wire na2273_2_i;
wire na2274_1;
wire na2274_1_i;
wire na2275_2;
wire na2275_2_i;
wire na2276_1;
wire na2276_1_i;
wire na2277_2;
wire na2277_2_i;
wire na2278_1;
wire na2278_1_i;
wire na2279_2;
wire na2279_2_i;
wire na2280_1;
wire na2280_1_i;
wire na2281_2;
wire na2281_2_i;
wire na2282_1;
wire na2282_1_i;
wire na2283_2;
wire na2283_2_i;
wire na2284_1;
wire na2284_1_i;
wire na2285_2;
wire na2285_2_i;
wire na2286_1;
wire na2286_1_i;
wire na2287_2;
wire na2287_2_i;
wire na2288_1;
wire na2288_1_i;
wire na2289_1;
wire na2289_1_i;
wire na2290_1;
wire na2290_1_i;
wire na2355_2;
wire na2355_2_i;
wire na2356_1;
wire na2356_1_i;
wire na2357_2;
wire na2357_2_i;
wire na2358_1;
wire na2358_1_i;
wire na2359_2;
wire na2359_2_i;
wire na2360_1;
wire na2360_1_i;
wire na2361_2;
wire na2361_2_i;
wire na2362_1;
wire na2362_1_i;
wire na2363_2;
wire na2363_2_i;
wire na2364_1;
wire na2364_1_i;
wire na2365_2;
wire na2365_2_i;
wire na2366_1;
wire na2366_1_i;
wire na2367_2;
wire na2367_2_i;
wire na2368_1;
wire na2368_1_i;
wire na2369_2;
wire na2369_2_i;
wire na2370_1;
wire na2370_1_i;
wire na2371_2;
wire na2371_2_i;
wire na2372_1;
wire na2372_1_i;
wire na2373_2;
wire na2373_2_i;
wire na2374_1;
wire na2374_1_i;
wire na2375_2;
wire na2375_2_i;
wire na2376_1;
wire na2376_1_i;
wire na2377_2;
wire na2377_2_i;
wire na2378_1;
wire na2378_1_i;
wire na2379_2;
wire na2379_2_i;
wire na2380_1;
wire na2380_1_i;
wire na2381_2;
wire na2381_2_i;
wire na2382_1;
wire na2382_1_i;
wire na2383_2;
wire na2383_2_i;
wire na2384_1;
wire na2384_1_i;
wire na2385_2;
wire na2385_2_i;
wire na2386_1;
wire na2386_1_i;
wire na2402_2;
wire na2402_2_i;
wire na2403_1;
wire na2403_1_i;
wire na2404_2;
wire na2404_2_i;
wire na2405_1;
wire na2405_1_i;
wire na2406_2;
wire na2406_2_i;
wire na2407_1;
wire na2407_1_i;
wire na2408_2;
wire na2408_2_i;
wire na2409_1;
wire na2409_1_i;
wire na2410_2;
wire na2410_2_i;
wire na2411_1;
wire na2411_1_i;
wire na2412_2;
wire na2412_2_i;
wire na2413_1;
wire na2413_1_i;
wire na2414_2;
wire na2414_2_i;
wire na2415_1;
wire na2415_1_i;
wire na2416_2;
wire na2416_2_i;
wire na2417_1;
wire na2417_1_i;
wire na2418_2;
wire na2418_2_i;
wire na2419_1;
wire na2419_1_i;
wire na2420_2;
wire na2420_2_i;
wire na2421_1;
wire na2421_1_i;
wire na2422_2;
wire na2422_2_i;
wire na2423_1;
wire na2423_1_i;
wire na2424_2;
wire na2424_2_i;
wire na2425_1;
wire na2425_1_i;
wire na2426_2;
wire na2426_2_i;
wire na2427_1;
wire na2427_1_i;
wire na2428_2;
wire na2428_2_i;
wire na2429_2;
wire na2429_2_i;
wire na2430_2;
wire na2430_2_i;
wire na2431_1;
wire na2431_1_i;
wire na2432_2;
wire na2432_2_i;
wire na2433_1;
wire na2433_1_i;
wire na2918_2;
wire na2918_2_i;
wire na2919_1;
wire na2919_1_i;
wire na2920_2;
wire na2920_2_i;
wire na2921_1;
wire na2921_1_i;
wire na2922_2;
wire na2922_2_i;
wire na2923_1;
wire na2923_1_i;
wire na2924_2;
wire na2924_2_i;
wire na2925_1;
wire na2925_1_i;
wire na2926_2;
wire na2926_2_i;
wire na2927_1;
wire na2927_1_i;
wire na2928_2;
wire na2928_2_i;
wire na2929_1;
wire na2929_1_i;
wire na2930_2;
wire na2930_2_i;
wire na2931_1;
wire na2931_1_i;
wire na2932_2;
wire na2932_2_i;
wire na2933_1;
wire na2933_1_i;
wire na2934_2;
wire na2934_2_i;
wire na2935_1;
wire na2935_1_i;
wire na2936_2;
wire na2936_2_i;
wire na2937_1;
wire na2937_1_i;
wire na2938_2;
wire na2938_2_i;
wire na2939_1;
wire na2939_1_i;
wire na2940_2;
wire na2940_2_i;
wire na2941_1;
wire na2941_1_i;
wire na2942_2;
wire na2942_2_i;
wire na2943_1;
wire na2943_1_i;
wire na2944_2;
wire na2944_2_i;
wire na2945_1;
wire na2945_1_i;
wire na2946_2;
wire na2946_2_i;
wire na2947_1;
wire na2947_1_i;
wire na2948_2;
wire na2948_2_i;
wire na2949_1;
wire na2949_1_i;
wire na3142_2;
wire na3142_2_i;
wire na3143_1;
wire na3143_1_i;
wire na3144_2;
wire na3144_2_i;
wire na3145_1;
wire na3145_1_i;
wire na3154_2;
wire na3154_2_i;
wire na3155_1;
wire na3155_1_i;
wire na3156_2;
wire na3156_2_i;
wire na3157_1;
wire na3157_1_i;
wire na3158_2;
wire na3158_2_i;
wire na3159_1;
wire na3159_1_i;
wire na3160_2;
wire na3160_2_i;
wire na3161_1;
wire na3161_1_i;
wire na3165_2;
wire na3165_2_i;
wire na3166_1;
wire na3166_1_i;
wire na3167_2;
wire na3167_2_i;
wire na3168_1;
wire na3168_1_i;
wire na3169_2;
wire na3169_2_i;
wire na3170_1;
wire na3170_1_i;
wire na3171_2;
wire na3171_2_i;
wire na3172_1;
wire na3172_1_i;
wire na3173_2;
wire na3173_2_i;
wire na3174_1;
wire na3174_1_i;
wire na3175_2;
wire na3175_2_i;
wire na3176_1;
wire na3176_1_i;
wire na3177_1;
wire na3177_1_i;
wire na3178_1;
wire na3178_1_i;
wire na3179_2;
wire na3179_2_i;
wire na3180_1;
wire na3180_1_i;
wire na3196_2;
wire na3196_2_i;
wire na3198_1;
wire na3198_1_i;
wire na3199_2;
wire na3199_2_i;
wire na3200_1;
wire na3200_1_i;
wire na3201_2;
wire na3201_2_i;
wire na3202_1;
wire na3202_1_i;
wire na3203_2;
wire na3203_2_i;
wire na3204_1;
wire na3204_1_i;
wire na3205_2;
wire na3205_2_i;
wire na3206_1;
wire na3206_1_i;
wire na3207_2;
wire na3207_2_i;
wire na3208_1;
wire na3208_1_i;
wire na3209_2;
wire na3209_2_i;
wire na3210_1;
wire na3210_1_i;
wire na3211_2;
wire na3211_2_i;
wire na3212_1;
wire na3212_1_i;
wire na3213_2;
wire na3213_2_i;
wire na3223_1;
wire na3223_1_i;
wire na3235_2;
wire na3235_2_i;
wire na3237_1;
wire na3237_1_i;
wire na3238_2;
wire na3238_2_i;
wire na3239_1;
wire na3239_1_i;
wire na3240_2;
wire na3240_2_i;
wire na3241_1;
wire na3241_1_i;
wire na3242_2;
wire na3242_2_i;
wire na3243_1;
wire na3243_1_i;
wire na3244_2;
wire na3244_2_i;
wire na3248_1;
wire na3249_1;
wire na3250_1;
wire na3251_1;
wire na3252_1;
wire na3253_1;
wire na3254_1;
wire na3255_1;
wire na3256_1;
wire na3257_1;
wire na3258_1;
wire na3259_1;
wire na3260_1;
wire na3261_1;
wire na3262_1;
wire na3263_1;
wire na3264_1;
wire na3265_1;
wire na3266_1;
wire na3267_1;
wire na3268_1;
wire na3269_1;
wire na3270_1;
wire na3271_1;
wire na3272_1;
wire na3273_1;
wire na3274_1;
wire na3275_1;
wire na3276_1;
wire na3277_1;
wire na3278_1;
wire na3279_1;
wire na3280_1;
wire na3281_1;
wire na3289_1;
wire na3290_1;
wire na3290_2;
wire na3292_2;
wire na3293_1;
wire na3294_2;
wire na3296_1;
wire na3296_4;
wire na3297_1;
wire na3298_1;
wire na3298_2;
wire na3300_1;
wire na3301_2;
wire na3303_1;
wire na3303_2;
wire na3305_2;
wire na3306_2;
wire na3308_1;
wire na3308_2;
wire na3310_1;
wire na3311_2;
wire na3313_1;
wire na3313_2;
wire na3315_1;
wire na3316_2;
wire na3318_1;
wire na3318_2;
wire na3320_1;
wire na3321_1;
wire na3323_1;
wire na3323_2;
wire na3325_1;
wire na3326_2;
wire na3328_1;
wire na3328_2;
wire na3330_1;
wire na3331_2;
wire na3333_1;
wire na3333_2;
wire na3335_2;
wire na3336_2;
wire na3338_1;
wire na3338_2;
wire na3340_2;
wire na3341_1;
wire na3343_1;
wire na3343_2;
wire na3345_2;
wire na3346_1;
wire na3348_1;
wire na3348_2;
wire na3350_1;
wire na3351_1;
wire na3353_1;
wire na3353_2;
wire na3355_2;
wire na3356_1;
wire na3358_1;
wire na3358_2;
wire na3360_2;
wire na3361_1;
wire na3363_1;
wire na3363_2;
wire na3365_2;
wire na3366_1;
wire na3368_1;
wire na3368_2;
wire na3370_1;
wire na3371_1;
wire na3373_1;
wire na3373_2;
wire na3375_2;
wire na3376_1;
wire na3378_1;
wire na3378_2;
wire na3380_2;
wire na3381_1;
wire na3383_1;
wire na3383_2;
wire na3385_2;
wire na3386_2;
wire na3388_1;
wire na3388_2;
wire na3390_2;
wire na3391_1;
wire na3393_1;
wire na3393_2;
wire na3395_2;
wire na3396_1;
wire na3398_1;
wire na3398_2;
wire na3400_2;
wire na3401_1;
wire na3403_1;
wire na3403_2;
wire na3405_1;
wire na3406_1;
wire na3408_1;
wire na3408_2;
wire na3410_2;
wire na3411_1;
wire na3413_1;
wire na3413_2;
wire na3415_2;
wire na3416_1;
wire na3418_1;
wire na3418_2;
wire na3420_2;
wire na3421_2;
wire na3423_1;
wire na3423_2;
wire na3425_1;
wire na3426_2;
wire na3428_1;
wire na3428_2;
wire na3430_1;
wire na3431_2;
wire na3433_1;
wire na3433_2;
wire na3435_1;
wire na3436_2;
wire na3438_1;
wire na3438_2;
wire na3440_1;
wire na3441_2;
wire na3443_1;
wire na3443_2;
wire na3445_1;
wire na3446_2;
wire na3448_1;
wire na3448_2;
wire na3450_2;
wire na3451_2;
wire na3453_1;
wire na3454_2;
wire na3456_1;
wire na3456_2;
wire na3457_1;
wire na3457_2;
wire na3459_1;
wire na3460_2;
wire na3463_1;
wire na3466_1;
wire na3467_1;
wire na3468_2;
wire na3469_1;
wire na3470_1;
wire na3470_2;
wire na3471_2;
wire na3472_1;
wire na3475_1;
wire na3475_2;
wire na3477_1;
wire na3477_2;
wire na3478_2;
wire na3480_2;
wire na3481_2;
wire na3485_1;
wire na3487_2;
wire na3489_1;
wire na3490_2;
wire na3494_1;
wire na3496_1;
wire na3497_2;
wire na3500_1;
wire na3501_1;
wire na3502_1;
wire na3504_2;
wire na3505_1;
wire na3509_2;
wire na3510_2;
wire na3515_1;
wire na3519_2;
wire na3520_1;
wire na3524_2;
wire na3526_2;
wire na3527_2;
wire na3530_1;
wire na3531_1;
wire na3531_2;
wire na3536_1;
wire na3536_2;
wire na3541_1;
wire na3543_2;
wire na3544_1;
wire na3544_2;
wire na3548_2;
wire na3550_2;
wire na3551_1;
wire na3551_2;
wire na3555_1;
wire na3555_2;
wire na3560_1;
wire na3561_1;
wire na3562_2;
wire na3563_1;
wire na3563_2;
wire na3569_1;
wire na3571_2;
wire na3572_1;
wire na3572_2;
wire na3576_1;
wire na3577_1;
wire na3579_1;
wire na3580_1;
wire na3580_2;
wire na3585_1;
wire na3586_1;
wire na3588_2;
wire na3589_1;
wire na3589_2;
wire na3594_1;
wire na3594_2;
wire na3599_1;
wire na3601_2;
wire na3602_1;
wire na3602_2;
wire na3606_1;
wire na3607_1;
wire na3608_2;
wire na3609_1;
wire na3609_2;
wire na3614_1;
wire na3619_1;
wire na3619_2;
wire na3621_1;
wire na3622_2;
wire na3624_1;
wire na3625_1;
wire na3625_2;
wire na3630_2;
wire na3632_1;
wire na3633_1;
wire na3633_2;
wire na3637_1;
wire na3638_2;
wire na3639_1;
wire na3640_1;
wire na3640_2;
wire na3646_1;
wire na3646_2;
wire na3651_1;
wire na3656_1;
wire na3656_2;
wire na3657_1;
wire na3659_2;
wire na3661_1;
wire na3662_1;
wire na3662_2;
wire na3666_2;
wire na3668_2;
wire na3669_1;
wire na3669_2;
wire na3673_1;
wire na3673_2;
wire na3675_1;
wire na3679_1;
wire na3680_2;
wire na3681_1;
wire na3682_1;
wire na3682_2;
wire na3688_2;
wire na3690_1;
wire na3691_1;
wire na3691_2;
wire na3695_1;
wire na3695_2;
wire na3700_2;
wire na3701_1;
wire na3702_1;
wire na3705_1;
wire na3705_2;
wire na3706_1;
wire na3711_1;
wire na3711_2;
wire na3715_1;
wire na3716_2;
wire na3717_1;
wire na3718_2;
wire na3719_1;
wire na3720_2;
wire na3721_1;
wire na3722_2;
wire na3723_1;
wire na3723_2;
wire na3724_1;
wire na3728_1;
wire na3728_2;
wire na3729_2;
wire na3730_1;
wire na3732_2;
wire na3734_1;
wire na3735_1;
wire na3736_1;
wire na3737_2;
wire na3738_1;
wire na3739_2;
wire na3740_1;
wire na3741_2;
wire na3742_2;
wire na3743_2;
wire na3744_1;
wire na3744_2;
wire na3745_1;
wire na3750_2;
wire na3752_1;
wire na3753_1;
wire na3753_2;
wire na3756_2;
wire na3757_1;
wire na3758_1;
wire na3759_1;
wire na3759_2;
wire na3763_1;
wire na3763_2;
wire na3765_1;
wire na3765_2;
wire na3766_1;
wire na3766_2;
wire na3767_1;
wire na3768_1;
wire na3768_2;
wire na3769_2;
wire na3770_1;
wire na3771_2;
wire na3772_1;
wire na3774_2;
wire na3775_1;
wire na3776_2;
wire na3777_1;
wire na3778_2;
wire na3779_1;
wire na3780_2;
wire na3781_2;
wire na3782_2;
wire na3783_1;
wire na3786_2;
wire na3790_1;
wire na3792_2;
wire na3793_1;
wire na3793_2;
wire na3796_1;
wire na3798_1;
wire na3800_1;
wire na3800_2;
wire na3801_1;
wire na3802_2;
wire na3804_1;
wire na3806_2;
wire na3808_1;
wire na3809_2;
wire na3811_2;
wire na3813_2;
wire na3814_1;
wire na3815_2;
wire na3816_1;
wire na3817_2;
wire na3818_1;
wire na3819_1;
wire na3820_1;
wire na3821_1;
wire na3822_2;
wire na3871_1;
wire na3871_2;
wire na3872_1;
wire na3873_2;
wire na3874_1;
wire na3875_2;
wire na3876_2;
wire na3877_1;
wire na3878_2;
wire na3952_1;
wire na3953_2;
wire na3954_1;
wire na3955_2;
wire na3956_2;
wire na3958_1;
wire na3959_1;
wire na3960_2;
wire na3961_1;
wire na3962_2;
wire na3963_1;
wire na3964_2;
wire na3965_1;
wire na3966_1;
wire na3967_1;
wire na3967_2;
wire na3968_1;
wire na3970_1;
wire na3971_1;
wire na3972_1;
wire na3973_2;
wire na3974_2;
wire na3975_2;
wire na3976_1;
wire na3977_2;
wire na3983_1;
wire na3984_2;
wire na3985_1;
wire na3986_1;
wire na3987_2;
wire na3988_1;
wire na3989_2;
wire na3990_1;
wire na3991_2;
wire na3994_1;
wire na3995_1;
wire na3996_2;
wire na3997_1;
wire na3998_2;
wire na3999_2;
wire na4000_2;
wire na4001_2;
wire na4003_2;
wire na4005_2;
wire na4006_1;
wire na4006_2;
wire na4013_1;
wire na4014_1;
wire na4015_1;
wire na4016_2;
wire na4025_1;
wire na4025_2;
wire na4026_1;
wire na4028_2;
wire na4029_1;
wire na4030_1;
wire na4031_1;
wire na4032_2;
wire na4033_1;
wire na4034_2;
wire na4035_2;
wire na4041_1;
wire na4041_2;
wire na4042_2;
wire na4044_2;
wire na4045_1;
wire na4046_2;
wire na4047_1;
wire na4048_2;
wire na4057_1;
wire na4057_2;
wire na4058_2;
wire na4060_1;
wire na4061_1;
wire na4063_2;
wire na4065_1;
wire na4066_1;
wire na4066_2;
wire na4072_1;
wire na4072_2;
wire na4073_2;
wire na4075_1;
wire na4076_2;
wire na4077_1;
wire na4078_2;
wire na4081_2;
wire na4084_2;
wire na4088_2;
wire na4089_1;
wire na4091_1;
wire na4093_1;
wire na4103_2;
wire na4104_1;
wire na4105_2;
wire na4106_1;
wire na4106_2;
wire na4108_1;
wire na4109_2;
wire na4112_1;
wire na4114_1;
wire na4115_1;
wire na4116_2;
wire na4117_1;
wire na4119_1;
wire na4120_1;
wire na4121_2;
wire na4122_1;
wire na4124_1;
wire na4125_1;
wire na4126_1;
wire na4127_1;
wire na4129_2;
wire na4130_1;
wire na4131_1;
wire na4133_1;
wire na4134_1;
wire na4138_1;
wire na4142_2;
wire na4143_1;
wire na4143_2;
wire na4148_1;
wire na4154_1;
wire na4155_1;
wire na4156_1;
wire na4157_2;
wire na4158_2;
wire na4159_2;
wire na4160_2;
wire na4161_2;
wire na4162_2;
wire na4163_2;
wire na4164_2;
wire na4165_2;
wire na4166_2;
wire na4167_2;
wire na4168_2;
wire na4169_2;
wire na4170_2;
wire na4171_2;
wire na4172_2;
wire na4173_2;
wire na4174_2;
wire na4175_2;
wire na4176_2;
wire na4177_2;
wire na4178_2;
wire na4179_2;
wire na4180_2;
wire na4181_2;
wire na4182_2;
wire na4183_2;
wire na4184_2;
wire na4185_2;
wire na4186_2;
wire na4187_2;
wire na4188_2;
wire na4189_2;
wire na4190_2;
wire na4191_2;
wire na4192_2;
wire na4193_2;
wire na4194_2;
wire na4195_2;
wire na4196_2;
wire na4197_2;
wire na4198_2;
wire na4199_2;
wire na4200_2;
wire na4201_2;
wire na4202_2;
wire na4203_2;
wire na4204_2;
wire na4205_2;
wire na4206_2;
wire na4207_2;
wire na4208_2;
wire na4209_2;
wire na4210_2;
wire na4211_2;
wire na4212_2;
wire na4213_2;
wire na4214_2;
wire na4215_2;
wire na4216_2;
wire na4217_2;
wire na4218_2;
wire na4219_2;
wire na4220_2;
wire na4221_2;
wire na4222_2;
wire na4223_2;
wire na4224_2;
wire na4225_2;
wire na4226_2;
wire na4227_2;
wire na4228_2;
wire na4229_2;
wire na4230_2;
wire na4231_2;
wire na4232_2;
wire na4233_2;
wire na4234_2;
wire na4235_2;
wire na4236_2;
wire na4237_2;
wire na4238_2;
wire na4239_2;
wire na4240_2;
wire na4241_2;
wire na4242_2;
wire na4243_2;
wire na4244_2;
wire na4245_2;
wire na4246_2;
wire na4247_2;
wire na4248_2;
wire na4249_2;
wire na4250_2;
wire na4251_2;
wire na4252_2;
wire na4253_2;
wire na4254_2;
wire na4255_2;
wire na4256_2;
wire na4257_2;
wire na4258_2;
wire na4259_2;
wire na4260_2;
wire na4261_2;
wire na4262_2;
wire na4263_2;
wire na4264_2;
wire na4265_2;
wire na4266_2;
wire na4267_2;
wire na4268_2;
wire na4269_2;
wire na4270_2;
wire na4271_2;
wire na4272_2;
wire na4273_2;
wire na4274_2;
wire na4275_2;
wire na4276_2;
wire na4277_2;
wire na4278_2;
wire na4279_2;
wire na4280_2;
wire na4281_2;
wire na4282_2;
wire na4283_2;
wire na4284_2;
wire na4285_2;
wire na4286_2;
wire na4287_2;
wire na4288_2;
wire na4289_2;
wire na4290_2;
wire na4291_2;
wire na4292_2;
wire na4293_2;
wire na4294_2;
wire na4295_2;
wire na4296_2;
wire na4297_2;
wire na4298_2;
wire na4299_2;
wire na4300_2;
wire na4301_2;
wire na4302_2;
wire na4303_2;
wire na4304_2;
wire na4305_2;
wire na4306_2;
wire na4307_2;
wire na4308_2;
wire na4309_2;
wire na4310_2;
wire na4311_2;
wire na4312_2;
wire na4313_2;
wire na4314_2;
wire na4315_2;
wire na4316_2;
wire na4317_2;
wire na4318_2;
wire na4319_2;
wire na4320_2;
wire na4321_2;
wire na4322_2;
wire na4323_2;
wire na4324_2;
wire na4325_2;
wire na4326_2;
wire na4327_2;
wire na4328_2;
wire na4329_2;
wire na4330_2;
wire na4331_2;
wire na4332_2;
wire na4333_2;
wire na4334_2;
wire na4335_2;
wire na4336_2;
wire na4337_2;
wire na4338_2;
wire na4339_2;
wire na4340_2;
wire na4341_2;
wire na4342_2;
wire na4343_2;
wire na4344_2;
wire na4345_2;
wire na4346_2;
wire na4347_2;
wire na4348_2;
wire na4349_2;
wire na4350_2;
wire na4351_2;
wire na4352_2;
wire na4353_2;
wire na4354_2;
wire na4355_2;
wire na4356_2;
wire na4357_2;
wire na4358_2;
wire na4359_2;
wire na4360_2;
wire na4361_2;
wire na4362_2;
wire na4363_2;
wire na4364_2;
wire na4365_2;
wire na4366_2;
wire na4367_2;
wire na4368_2;
wire na4369_2;
wire na4370_2;
wire na4371_2;
wire na4372_2;
wire na4373_2;
wire na4374_2;
wire na4375_2;
wire na4376_2;
wire na4377_2;
wire na4378_2;
wire na4379_2;
wire na4380_2;
wire na4381_2;
wire na4382_2;
wire na4383_2;
wire na4384_2;
wire na4385_2;
wire na4386_2;
wire na4387_2;
wire na4388_2;
wire na4389_2;
wire na4390_2;
wire na4391_2;
wire na4392_2;
wire na4393_2;
wire na4394_2;
wire na4395_2;
wire na4396_2;
wire na4397_2;
wire na4398_2;
wire na4399_2;
wire na4400_2;
wire na4401_2;
wire na4402_2;
wire na4403_2;
wire na4404_2;
wire na4405_2;
wire na4406_2;
wire na4407_2;
wire na4408_2;
wire na4409_2;
wire na4410_2;
wire na4411_2;
wire na4412_2;
wire na4413_2;
wire na4414_2;
wire na4415_2;
wire na4416_2;
wire na4417_2;
wire na4418_2;
wire na4419_2;
wire na4420_2;
wire na4421_2;
wire na4422_2;
wire na4423_2;
wire na4424_2;
wire na4425_2;
wire na4426_2;
wire na4427_2;
wire na4428_2;
wire na4429_2;
wire na4430_2;
wire na4431_2;
wire na4432_2;
wire na4433_2;
wire na4512_1;
wire na4512_2;
wire na4512_3;
wire na4512_6;
wire na4158_10;
wire na4159_10;
wire na4160_10;
wire na4161_10;
wire na4162_10;
wire na4163_10;
wire na4164_10;

CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a1 ( .PCLK0(na1_1), .PCLK1(_d0), .PCLK2(_d1), .PCLK3(_d2), .CLK0(na3280_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0), .SER_CLK(1'b0),
                 .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_AND/D///      x86y83     80'h40_E400_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1337_1), .IN7(na1872_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2_2 ( .OUT(na2_1), .CLK(1'b0), .EN(~na1467_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                   .D_IN(na2_1_i) );
// C_AND/D//AND/D      x81y83     80'h40_E400_80_0000_0C88_ACF4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3_1 ( .OUT(na3_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1337_1), .IN7(na1872_2), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3_2 ( .OUT(na3_1), .CLK(1'b0), .EN(~na1467_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                   .D_IN(na3_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3_4 ( .OUT(na3_2_i), .IN1(~na3_2), .IN2(na1337_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3_5 ( .OUT(na3_2), .CLK(1'b0), .EN(~na1467_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                   .D_IN(na3_2_i) );
// C_AND/D//AND/D      x85y88     80'h40_E400_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1337_1), .IN7(1'b1), .IN8(na1874_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a5_2 ( .OUT(na5_1), .CLK(1'b0), .EN(~na1467_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                   .D_IN(na5_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2_i), .IN1(1'b1), .IN2(na1337_1), .IN3(1'b1), .IN4(na1874_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a5_5 ( .OUT(na5_2), .CLK(1'b0), .EN(~na1467_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                   .D_IN(na5_2_i) );
// C_AND/D///      x91y91     80'h40_E400_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1337_1), .IN7(na1876_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a6_2 ( .OUT(na6_1), .CLK(1'b0), .EN(~na1467_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                   .D_IN(na6_1_i) );
// C_AND////      x154y66     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na539_1), .IN6(1'b1), .IN7(1'b1), .IN8(na549_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x156y66     80'h40_E800_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2_i), .IN1(na1878_1), .IN2(1'b1), .IN3(1'b1), .IN4(na7_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a9_5 ( .OUT(na9_2), .CLK(1'b0), .EN(na1468_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                   .D_IN(na9_2_i) );
// C_AND/D//AND/D      x153y71     80'h40_E800_80_0000_0C88_CAC5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1878_2), .IN6(1'b1), .IN7(1'b1), .IN8(na7_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a10_2 ( .OUT(na10_1), .CLK(1'b0), .EN(na1468_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na10_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a10_4 ( .OUT(na10_2_i), .IN1(~na10_2), .IN2(1'b1), .IN3(1'b1), .IN4(na7_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a10_5 ( .OUT(na10_2), .CLK(1'b0), .EN(na1468_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na10_2_i) );
// C_AND/D//AND/D      x153y74     80'h40_E800_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1880_2), .IN7(1'b1), .IN8(na7_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a12_2 ( .OUT(na12_1), .CLK(1'b0), .EN(na1468_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na12_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a12_4 ( .OUT(na12_2_i), .IN1(1'b1), .IN2(na1880_1), .IN3(1'b1), .IN4(na7_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a12_5 ( .OUT(na12_2), .CLK(1'b0), .EN(na1468_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na12_2_i) );
// C_OR/D///      x98y88     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1_i), .IN1(na14_1), .IN2(na24_1), .IN3(na22_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3290_2), .IN8(na4369_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a13_2 ( .OUT(na13_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na13_1_i) );
// C_ORAND////      x107y73     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3292_2), .IN8(~na17_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y65     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a15_4 ( .OUT(na15_2), .IN1(~na16_2), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x109y67     80'h00_0060_00_0000_0C08_FF31
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a16_4 ( .OUT(na16_2), .IN1(~na1335_2), .IN2(~na4341_2), .IN3(1'b1), .IN4(~na1336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y80     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3293_1), .IN6(~na712_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x127y77     80'h00_0078_00_0000_0C88_C1F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a21_1 ( .OUT(na21_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1331_1), .IN6(~na1859_1), .IN7(1'b1), .IN8(na1332_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a21_4 ( .OUT(na21_2), .IN1(~na3294_2), .IN2(~na1859_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y83     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na648_1), .IN6(na744_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y86     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na592_1), .IN6(na551_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x116y78     80'h00_0078_00_0000_0CEE_3DCD
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1331_1), .IN6(na1859_1), .IN7(1'b0), .IN8(~na1332_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a25_4 ( .OUT(na25_2), .IN1(~na1331_1), .IN2(na1859_1), .IN3(1'b0), .IN4(na1332_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x131y81     80'h00_0078_00_0000_0C88_F8F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_1 ( .OUT(na26_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na21_1), .IN6(na1333_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a26_4 ( .OUT(na26_2), .IN1(na21_1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x124y81     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1_i), .IN1(na32_1), .IN2(na28_1), .IN3(na33_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3298_2), .IN8(na4370_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a27_2 ( .OUT(na27_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na27_1_i) );
// C_ORAND////      x127y80     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3300_1), .IN8(~na30_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y76     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3301_2), .IN6(~na713_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y81     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na553_1), .IN6(na593_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y77     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na745_1), .IN8(na649_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x133y95     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_1 ( .OUT(na34_1_i), .IN1(na39_1), .IN2(na35_2), .IN3(na3303_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3303_2),
                    .IN8(na38_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a34_2 ( .OUT(na34_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na34_1_i) );
// C_///ORAND/      x119y76     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a35_4 ( .OUT(na35_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na36_1), .IN4(na3305_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y83     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3306_2), .IN6(~na714_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y90     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na650_1), .IN8(na4231_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y85     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na594_1), .IN6(na554_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x127y63     80'h40_E800_00_0000_0EEE_E0EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a40_1 ( .OUT(na40_1_i), .IN1(na41_1), .IN2(1'b0), .IN3(na45_1), .IN4(na3308_2), .IN5(1'b0), .IN6(1'b0), .IN7(na44_1), .IN8(na3308_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a40_2 ( .OUT(na40_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na40_1_i) );
// C_ORAND////      x115y67     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3310_1), .IN8(~na42_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y60     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3311_2), .IN8(~na715_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y69     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na555_1), .IN6(na595_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y67     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na651_1), .IN6(na4232_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x108y68     80'h40_E800_00_0000_0EEE_CAEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1_i), .IN1(na3313_2), .IN2(1'b0), .IN3(na51_1), .IN4(na47_2), .IN5(na3313_1), .IN6(1'b0), .IN7(1'b0),
                    .IN8(na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a46_2 ( .OUT(na46_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na46_1_i) );
// C_///ORAND/      x110y66     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a47_4 ( .OUT(na47_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na48_1), .IN4(na3315_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y69     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3316_2), .IN8(~na716_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y70     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na652_1), .IN6(na748_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y73     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na556_1), .IN6(na596_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x94y70     80'h40_E800_00_0000_0EEE_AECA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a52_1 ( .OUT(na52_1_i), .IN1(na3318_2), .IN2(1'b0), .IN3(1'b0), .IN4(na53_1), .IN5(na3318_1), .IN6(na56_1), .IN7(na57_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a52_2 ( .OUT(na52_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na52_1_i) );
// C_ORAND////      x98y72     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3320_1), .IN8(~na54_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y72     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3321_1), .IN6(~na717_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y78     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a56_1 ( .OUT(na56_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na597_1), .IN6(na557_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x94y71     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na653_1), .IN6(na4233_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x105y63     80'h40_E800_00_0000_0EEE_AECA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1_i), .IN1(na3323_2), .IN2(1'b0), .IN3(1'b0), .IN4(na59_2), .IN5(na3323_1), .IN6(na62_1), .IN7(na63_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a58_2 ( .OUT(na58_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na58_1_i) );
// C_///ORAND/      x120y62     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a59_4 ( .OUT(na59_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na60_1), .IN4(na3325_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y63     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a60_1 ( .OUT(na60_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3326_2), .IN8(~na718_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y70     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na558_1), .IN6(na4222_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y65     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na4234_2), .IN8(na654_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x111y62     80'h40_E800_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1_i), .IN1(1'b0), .IN2(na65_1), .IN3(na69_1), .IN4(na3328_2), .IN5(1'b0), .IN6(1'b0), .IN7(na68_1), .IN8(na3328_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a64_2 ( .OUT(na64_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na64_1_i) );
// C_ORAND////      x119y64     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3330_1), .IN8(~na66_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y64     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3331_2), .IN8(~na719_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y65     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_1 ( .OUT(na68_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na751_1), .IN8(na655_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y67     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(1'b0), .IN7(na559_1), .IN8(na4224_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x104y81     80'h40_E800_00_0000_0EEE_CCAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1_i), .IN1(na71_2), .IN2(na3333_2), .IN3(na75_1), .IN4(1'b0), .IN5(1'b0), .IN6(na3333_1), .IN7(1'b0),
                    .IN8(na74_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a70_2 ( .OUT(na70_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na70_1_i) );
// C_///ORAND/      x99y77     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a71_4 ( .OUT(na71_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na72_1), .IN4(na3335_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y83     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_1 ( .OUT(na72_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na720_1), .IN6(~na3336_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y88     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na560_1), .IN6(na600_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y87     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na752_1), .IN8(na656_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x115y86     80'h40_E800_00_0000_0EEE_CCEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1_i), .IN1(1'b0), .IN2(na77_1), .IN3(na81_1), .IN4(na3338_2), .IN5(1'b0), .IN6(na80_1), .IN7(1'b0), .IN8(na3338_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a76_2 ( .OUT(na76_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na76_1_i) );
// C_ORAND////      x111y80     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a77_1 ( .OUT(na77_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na78_1), .IN8(na3340_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y85     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na721_1), .IN6(~na3341_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y88     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na561_1), .IN6(na601_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y87     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na753_1), .IN8(na657_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x110y88     80'h40_E800_00_0000_0EEE_CAEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a82_1 ( .OUT(na82_1_i), .IN1(1'b0), .IN2(na87_1), .IN3(na83_2), .IN4(na3343_2), .IN5(na86_1), .IN6(1'b0), .IN7(1'b0), .IN8(na3343_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a82_2 ( .OUT(na82_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na82_1_i) );
// C_///ORAND/      x106y77     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a83_4 ( .OUT(na83_2), .IN1(~na21_2), .IN2(1'b0), .IN3(na3345_2), .IN4(~na84_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y86     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3346_1), .IN6(~na722_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y87     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na602_1), .IN6(na562_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y88     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na754_1), .IN8(na4228_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x112y73     80'h40_E800_00_0000_0EEE_AECC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1_i), .IN1(1'b0), .IN2(na3348_2), .IN3(1'b0), .IN4(na89_1), .IN5(na92_1), .IN6(na3348_1), .IN7(na93_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a88_2 ( .OUT(na88_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na88_1_i) );
// C_ORAND////      x114y72     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na90_1), .IN8(na3350_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y73     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3351_1), .IN8(~na723_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y77     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na755_1), .IN6(na659_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y75     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na563_1), .IN6(na4225_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x105y73     80'h40_E800_00_0000_0EEE_0EAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1_i), .IN1(na95_2), .IN2(na3353_2), .IN3(na99_1), .IN4(1'b0), .IN5(na98_1), .IN6(na3353_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a94_2 ( .OUT(na94_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na94_1_i) );
// C_///ORAND/      x113y69     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a95_4 ( .OUT(na95_2), .IN1(~na21_2), .IN2(1'b0), .IN3(na3355_2), .IN4(~na96_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y74     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a96_1 ( .OUT(na96_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na724_1), .IN8(~na3356_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y79     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_1 ( .OUT(na98_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na564_1), .IN6(na604_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y81     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na756_1), .IN6(na660_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y70     80'h40_E800_00_0000_0EEE_CCAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1_i), .IN1(na105_1), .IN2(na3358_2), .IN3(na101_1), .IN4(1'b0), .IN5(1'b0), .IN6(na3358_1), .IN7(1'b0),
                     .IN8(na104_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a100_2 ( .OUT(na100_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na100_1_i) );
// C_ORAND////      x100y73     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a101_1 ( .OUT(na101_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na102_1), .IN8(na3360_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y75     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3361_1), .IN6(~na725_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y78     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na605_1), .IN6(na4204_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y77     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na757_1), .IN8(na661_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x96y68     80'h40_E800_00_0000_0EEE_ECE0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na4371_2), .IN4(na107_2), .IN5(1'b0), .IN6(na111_1), .IN7(na110_1),
                     .IN8(na3363_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a106_2 ( .OUT(na106_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na106_1_i) );
// C_///ORAND/      x98y66     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a107_4 ( .OUT(na107_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na108_1), .IN4(na3365_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y67     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_1 ( .OUT(na108_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na726_1), .IN6(~na3366_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x92y67     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na662_1), .IN6(na758_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y72     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na606_1), .IN6(na4205_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x102y64     80'h40_E800_00_0000_0EEE_ECCA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1_i), .IN1(na113_1), .IN2(1'b0), .IN3(1'b0), .IN4(na117_1), .IN5(1'b0), .IN6(na4372_2), .IN7(na116_1),
                     .IN8(na3368_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a112_2 ( .OUT(na112_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na112_1_i) );
// C_ORAND////      x101y65     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na114_1), .IN8(na3370_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y63     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a114_1 ( .OUT(na114_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3371_1), .IN6(~na727_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y65     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a116_1 ( .OUT(na116_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na663_1), .IN8(na759_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y70     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na4207_2), .IN6(na607_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x143y96     80'h40_E800_00_0000_0EEE_0EEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1_i), .IN1(na3373_2), .IN2(1'b0), .IN3(na123_1), .IN4(na119_2), .IN5(na3373_1), .IN6(na122_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a118_2 ( .OUT(na118_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na118_1_i) );
// C_///ORAND/      x138y88     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a119_4 ( .OUT(na119_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na120_1), .IN4(na3375_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y93     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a120_1 ( .OUT(na120_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na728_1), .IN8(~na3376_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y88     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na568_1), .IN6(na608_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y93     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na760_1), .IN6(na664_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x130y96     80'h40_E800_00_0000_0EEE_0EEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a124_1 ( .OUT(na124_1_i), .IN1(na3378_2), .IN2(1'b0), .IN3(na129_1), .IN4(na125_1), .IN5(na3378_1), .IN6(na128_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a124_2 ( .OUT(na124_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na124_1_i) );
// C_ORAND////      x132y92     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na126_1), .IN8(na3380_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y91     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a126_1 ( .OUT(na126_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3381_1), .IN6(~na729_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y96     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na569_1), .IN6(na609_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y95     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a129_1 ( .OUT(na129_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na665_1), .IN6(na4235_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x127y95     80'h40_E800_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a130_1 ( .OUT(na130_1_i), .IN1(1'b0), .IN2(na131_2), .IN3(na3383_2), .IN4(na135_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3383_1),
                     .IN8(na134_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a130_2 ( .OUT(na130_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na130_1_i) );
// C_///ORAND/      x133y88     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a131_4 ( .OUT(na131_2), .IN1(~na21_2), .IN2(1'b0), .IN3(na3385_2), .IN4(~na132_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y90     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a132_1 ( .OUT(na132_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3386_2), .IN8(~na730_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y94     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(1'b0), .IN7(na4209_2), .IN8(na610_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y94     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a135_1 ( .OUT(na135_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na4236_2), .IN8(na666_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x138y94     80'h40_E800_00_0000_0EEE_CCAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1_i), .IN1(na141_1), .IN2(na3388_2), .IN3(na137_1), .IN4(1'b0), .IN5(1'b0), .IN6(na3388_1), .IN7(1'b0),
                     .IN8(na140_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a136_2 ( .OUT(na136_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na136_1_i) );
// C_ORAND////      x142y85     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a137_1 ( .OUT(na137_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na138_1), .IN8(na3390_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x136y91     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3391_1), .IN6(~na731_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y94     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na667_1), .IN8(na763_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y91     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na571_1), .IN6(na611_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x130y91     80'h40_E800_00_0000_0EEE_ACCE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a142_1 ( .OUT(na142_1_i), .IN1(na143_2), .IN2(na3393_2), .IN3(1'b0), .IN4(na147_1), .IN5(1'b0), .IN6(na3393_1), .IN7(na146_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a142_2 ( .OUT(na142_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na142_1_i) );
// C_///ORAND/      x125y85     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a143_4 ( .OUT(na143_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na144_1), .IN4(na3395_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y85     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a144_1 ( .OUT(na144_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3396_1), .IN6(~na732_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y85     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na572_1), .IN6(na612_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y88     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a147_1 ( .OUT(na147_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na668_1), .IN8(na764_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x128y87     80'h40_E800_00_0000_0EEE_ACAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1_i), .IN1(na149_1), .IN2(na3398_2), .IN3(na153_1), .IN4(1'b0), .IN5(1'b0), .IN6(na3398_1), .IN7(na152_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a148_2 ( .OUT(na148_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na148_1_i) );
// C_ORAND////      x123y81     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a149_1 ( .OUT(na149_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3400_2), .IN8(~na150_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x120y82     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3401_1), .IN6(~na733_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y83     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na613_1), .IN6(na573_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y87     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a153_1 ( .OUT(na153_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na765_1), .IN6(na669_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x110y64     80'h40_E800_00_0000_0EEE_CCAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1_i), .IN1(na159_1), .IN2(na3403_2), .IN3(na155_2), .IN4(1'b0), .IN5(1'b0), .IN6(na3403_1), .IN7(1'b0),
                     .IN8(na158_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a154_2 ( .OUT(na154_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na154_1_i) );
// C_///ORAND/      x118y67     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a155_4 ( .OUT(na155_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na156_1), .IN4(na3405_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y67     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a156_1 ( .OUT(na156_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3406_1), .IN8(~na734_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y70     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a158_1 ( .OUT(na158_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na614_1), .IN6(na4211_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y67     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a159_1 ( .OUT(na159_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na670_1), .IN6(na766_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x131y67     80'h40_E800_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_1 ( .OUT(na160_1_i), .IN1(1'b0), .IN2(na161_1), .IN3(na165_1), .IN4(na3408_2), .IN5(1'b0), .IN6(1'b0), .IN7(na164_1),
                     .IN8(na3408_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a160_2 ( .OUT(na160_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na160_1_i) );
// C_ORAND////      x125y68     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3410_2), .IN8(~na162_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x124y68     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a162_1 ( .OUT(na162_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3411_1), .IN8(~na735_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y69     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na575_1), .IN6(na4227_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y75     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_1 ( .OUT(na165_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na767_1), .IN6(na671_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x116y92     80'h40_E800_00_0000_0EEE_AACE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1_i), .IN1(na3413_2), .IN2(na167_2), .IN3(1'b0), .IN4(na171_1), .IN5(na3413_1), .IN6(1'b0), .IN7(na170_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a166_2 ( .OUT(na166_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na166_1_i) );
// C_///ORAND/      x115y84     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a167_4 ( .OUT(na167_2), .IN1(~na21_2), .IN2(1'b0), .IN3(na3415_2), .IN4(~na168_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y86     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3416_1), .IN8(~na736_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y87     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_1 ( .OUT(na170_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na584_1), .IN6(na4213_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y90     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a171_1 ( .OUT(na171_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na768_1), .IN8(na672_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x120y94     80'h40_E800_00_0000_0EEE_EACC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a172_1 ( .OUT(na172_1_i), .IN1(1'b0), .IN2(na173_1), .IN3(1'b0), .IN4(na3418_2), .IN5(na177_1), .IN6(1'b0), .IN7(na176_1),
                     .IN8(na3418_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a172_2 ( .OUT(na172_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na172_1_i) );
// C_ORAND////      x115y84     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na174_1), .IN8(na3420_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y87     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a174_1 ( .OUT(na174_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3421_2), .IN6(~na737_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y89     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a176_1 ( .OUT(na176_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na4214_2), .IN6(na585_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y91     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na4237_2), .IN6(na673_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x131y96     80'h40_E800_00_0000_0EEE_AAAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1_i), .IN1(na3423_2), .IN2(na179_2), .IN3(na183_1), .IN4(1'b0), .IN5(na3423_1), .IN6(1'b0), .IN7(na182_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a178_2 ( .OUT(na178_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na178_1_i) );
// C_///ORAND/      x125y86     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a179_4 ( .OUT(na179_2), .IN1(~na21_2), .IN2(1'b0), .IN3(na3425_1), .IN4(~na180_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y90     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3426_2), .IN6(~na738_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y91     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na586_1), .IN6(na4215_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y101     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na770_1), .IN8(na4229_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x114y83     80'h40_E800_00_0000_0EEE_ECCA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a184_1 ( .OUT(na184_1_i), .IN1(na185_1), .IN2(1'b0), .IN3(1'b0), .IN4(na3428_2), .IN5(1'b0), .IN6(na189_1), .IN7(na188_1),
                     .IN8(na3428_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a184_2 ( .OUT(na184_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na184_1_i) );
// C_ORAND////      x111y79     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a185_1 ( .OUT(na185_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na186_1), .IN8(na3430_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y83     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na739_1), .IN6(~na3431_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y85     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na579_1), .IN6(na587_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y86     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a189_1 ( .OUT(na189_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na4238_2), .IN6(na675_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x109y88     80'h40_E800_00_0000_0EEE_AACE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a190_1 ( .OUT(na190_1_i), .IN1(na3433_2), .IN2(na191_2), .IN3(1'b0), .IN4(na195_1), .IN5(na3433_1), .IN6(1'b0), .IN7(na194_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a190_2 ( .OUT(na190_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na190_1_i) );
// C_///ORAND/      x109y80     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a191_4 ( .OUT(na191_2), .IN1(~na21_2), .IN2(1'b0), .IN3(na3435_1), .IN4(~na192_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y86     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a192_1 ( .OUT(na192_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3436_2), .IN6(~na740_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y83     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(1'b0), .IN7(na4216_2), .IN8(na588_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y86     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a195_1 ( .OUT(na195_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na772_1), .IN6(na676_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x102y83     80'h40_E800_00_0000_0EEE_AECA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a196_1 ( .OUT(na196_1_i), .IN1(na3438_2), .IN2(1'b0), .IN3(1'b0), .IN4(na197_1), .IN5(na3438_1), .IN6(na201_1), .IN7(na200_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a196_2 ( .OUT(na196_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na196_1_i) );
// C_ORAND////      x104y80     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a197_1 ( .OUT(na197_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(~na198_1), .IN8(na3440_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y83     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a198_1 ( .OUT(na198_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3441_2), .IN6(~na741_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y87     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a200_1 ( .OUT(na200_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na589_1), .IN6(na4217_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y90     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a201_1 ( .OUT(na201_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na773_1), .IN6(na4230_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x103y71     80'h40_E800_00_0000_0EEE_AACE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1_i), .IN1(na3443_2), .IN2(na203_2), .IN3(1'b0), .IN4(na207_1), .IN5(na3443_1), .IN6(1'b0), .IN7(na206_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a202_2 ( .OUT(na202_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na202_1_i) );
// C_///ORAND/      x111y70     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a203_4 ( .OUT(na203_2), .IN1(~na21_2), .IN2(1'b0), .IN3(~na204_1), .IN4(na3445_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y69     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a204_1 ( .OUT(na204_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na742_1), .IN6(~na3446_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y75     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a206_1 ( .OUT(na206_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(na4218_2), .IN6(na590_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y76     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na678_1), .IN6(na774_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x105y68     80'h40_E800_00_0000_0EEE_0EEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_1 ( .OUT(na208_1_i), .IN1(na3448_2), .IN2(1'b0), .IN3(na209_1), .IN4(na213_1), .IN5(na3448_1), .IN6(na212_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a208_2 ( .OUT(na208_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na208_1_i) );
// C_ORAND////      x112y67     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a209_1 ( .OUT(na209_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_2), .IN6(1'b0), .IN7(na3450_2), .IN8(~na210_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x106y68     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a210_1 ( .OUT(na210_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3451_2), .IN6(~na743_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y72     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na679_1), .IN6(na775_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y72     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a213_1 ( .OUT(na213_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(1'b0), .IN7(na583_1), .IN8(na591_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x102y77     80'h40_E818_00_0000_0666_0AA3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1), .IN1(1'b0), .IN2(~na259_1), .IN3(na260_1), .IN4(1'b0), .IN5(na215_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a214_5 ( .OUT(na214_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na214_1) );
// C_XOR///XOR/      x87y71     80'h00_0078_00_0000_0C66_6C99
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a215_1 ( .OUT(na215_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na255_1), .IN7(na216_1), .IN8(na249_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a215_4 ( .OUT(na215_2), .IN1(na268_1), .IN2(~na291_1), .IN3(~na290_1), .IN4(na269_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y69     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a216_1 ( .OUT(na216_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na243_1), .IN8(na217_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y68     80'h00_0018_00_0040_0A72_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a217_1 ( .OUT(na217_1), .IN1(1'b1), .IN2(na4179_2), .IN3(1'b1), .IN4(na4185_2), .IN5(na3453_1), .IN6(~na241_1), .IN7(na240_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y80     80'h00_0018_00_0040_0AF9_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1), .IN1(na1811_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na228_1), .IN5(~na4373_2), .IN6(na1814_1), .IN7(na3454_2),
                     .IN8(~na4184_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x82y98     80'h00_0018_00_0040_0AE6_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a221_1 ( .OUT(na221_1), .IN1(1'b1), .IN2(~na4374_2), .IN3(~na225_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na223_2), .IN7(~na225_1),
                     .IN8(na3456_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x81y96     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a223_4 ( .OUT(na223_2), .IN1(~na1154_1), .IN2(na1166_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x86y93     80'h00_0078_00_0000_0C66_3A96
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_1 ( .OUT(na225_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1154_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1156_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a225_4 ( .OUT(na225_2), .IN1(na1154_1), .IN2(na1166_1), .IN3(na1160_1), .IN4(~na1164_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x85y94     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1154_1), .IN6(~na1166_1), .IN7(na1160_1),
                     .IN8(na1156_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x80y84     80'h00_0018_00_0000_0666_CA56
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a228_1 ( .OUT(na228_1), .IN1(na3459_1), .IN2(na223_2), .IN3(~na3460_2), .IN4(1'b0), .IN5(na229_1), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na231_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x87y97     80'h00_0018_00_0040_0C23_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(na3457_1), .IN2(~na4375_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3457_2), .IN6(1'b1), .IN7(na225_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x88y98     80'h00_0018_00_0040_0C26_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1), .IN1(1'b0), .IN2(~na1166_1), .IN3(na4320_2), .IN4(1'b0), .IN5(na1162_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na1156_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y97     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a233_4 ( .OUT(na233_2), .IN1(~na3470_2), .IN2(1'b1), .IN3(~na225_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x81y95     80'h00_0018_00_0000_0666_EA5D
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_1 ( .OUT(na234_1), .IN1(na3463_1), .IN2(~na223_2), .IN3(na236_1), .IN4(1'b1), .IN5(~na238_1), .IN6(1'b1), .IN7(~na4376_2),
                     .IN8(~na3456_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y97     80'h00_0018_00_0040_0A32_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_1 ( .OUT(na236_1), .IN1(~na3470_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3457_1), .IN6(~na4377_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y95     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_1 ( .OUT(na238_1), .IN1(1'b1), .IN2(na4432_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4318_2), .IN8(~na1156_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y78     80'h00_0018_00_0040_0AF1_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(~na234_1), .IN2(1'b1), .IN3(1'b1), .IN4(na228_1), .IN5(~na1811_1), .IN6(na1814_1), .IN7(na4360_2),
                     .IN8(na3466_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x80y73     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a240_4 ( .OUT(na240_2), .IN1(1'b0), .IN2(na223_2), .IN3(1'b0), .IN4(~na4106_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y74     80'h00_0018_00_0000_0C66_5C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_1 ( .OUT(na241_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na227_1), .IN7(~na242_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x86y89     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a242_4 ( .OUT(na242_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1158_1), .IN4(na1156_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y71     80'h00_0018_00_0040_0ABD_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1), .IN1(na244_1), .IN2(1'b1), .IN3(1'b1), .IN4(na245_1), .IN5(~na246_1), .IN6(na3467_1), .IN7(1'b1),
                     .IN8(~na248_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y89     80'h00_0018_00_0040_0AF4_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a244_1 ( .OUT(na244_1), .IN1(1'b1), .IN2(na1814_1), .IN3(1'b1), .IN4(~na228_1), .IN5(na1811_1), .IN6(na4182_2), .IN7(~na4183_2),
                     .IN8(na3468_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y76     80'h00_0018_00_0040_0AFC_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a245_1 ( .OUT(na245_1), .IN1(1'b1), .IN2(na1814_1), .IN3(na4183_2), .IN4(1'b1), .IN5(na1811_1), .IN6(na3469_1), .IN7(~na4360_2),
                     .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y85     80'h00_0018_00_0000_0C66_3C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_1 ( .OUT(na246_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1151_1), .IN7(1'b0), .IN8(~na4380_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x80y82     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a248_4 ( .OUT(na248_2), .IN1(1'b0), .IN2(1'b0), .IN3(na225_1), .IN4(na4181_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x82y72     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a249_4 ( .OUT(na249_2), .IN1(~na252_1), .IN2(na251_1), .IN3(na254_1), .IN4(na250_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x82y88     80'h00_0018_00_0040_0AD3_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a250_1 ( .OUT(na250_1), .IN1(na3470_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_1), .IN5(~na244_1), .IN6(1'b1), .IN7(na4378_2),
                     .IN8(na3456_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y86     80'h00_0018_00_0040_0A7A_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a251_1 ( .OUT(na251_1), .IN1(1'b1), .IN2(na239_1), .IN3(1'b1), .IN4(na245_1), .IN5(na3471_2), .IN6(~na4432_2), .IN7(na225_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y85     80'h00_0018_00_0040_0ABD_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1), .IN1(na244_1), .IN2(1'b1), .IN3(1'b1), .IN4(na245_1), .IN5(~na4187_2), .IN6(na3472_1), .IN7(1'b1),
                     .IN8(~na253_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y92     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a253_1 ( .OUT(na253_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3470_2), .IN6(1'b0), .IN7(1'b0), .IN8(na3456_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x86y85     80'h00_0018_00_0040_0AE9_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(1'b1), .IN2(~na239_1), .IN3(1'b1), .IN4(~na218_1), .IN5(1'b1), .IN6(na4379_2), .IN7(na225_2),
                     .IN8(~na4106_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x85y86     80'h00_0018_00_0000_0666_EFA7
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a255_1 ( .OUT(na255_1), .IN1(na244_1), .IN2(na4432_2), .IN3(~na256_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na225_2),
                     .IN8(~na245_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x82y89     80'h00_0018_00_0040_0ABC_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1), .IN1(1'b1), .IN2(~na239_1), .IN3(1'b1), .IN4(na218_1), .IN5(na3470_2), .IN6(na4374_2), .IN7(1'b1),
                     .IN8(~na253_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y88     80'h00_0018_00_0040_0ABD_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a259_1 ( .OUT(na259_1), .IN1(1'b1), .IN2(~na4179_2), .IN3(1'b1), .IN4(na4380_2), .IN5(~na244_1), .IN6(na3477_1), .IN7(1'b1),
                     .IN8(~na4317_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x84y83     80'h00_0018_00_0040_0A7E_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1), .IN1(1'b1), .IN2(na4188_2), .IN3(1'b1), .IN4(na4185_2), .IN5(na3478_2), .IN6(~na4189_2), .IN7(~na240_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x127y72     80'h00_0060_00_0000_0C08_FF3D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a261_4 ( .OUT(na261_2), .IN1(~na262_1), .IN2(na3480_2), .IN3(1'b0), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y75     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3481_2), .IN8(~na1133_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x121y76     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a263_1 ( .OUT(na263_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_1), .IN6(~na2051_2), .IN7(~na2019_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x115y77     80'h40_E818_00_0000_0666_C3A0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a264_1 ( .OUT(na264_1), .IN1(1'b0), .IN2(1'b0), .IN3(na273_1), .IN4(1'b0), .IN5(1'b0), .IN6(~na255_1), .IN7(1'b0), .IN8(na265_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a264_5 ( .OUT(na264_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na264_1) );
// C_XOR////      x84y80     80'h00_0018_00_0000_0666_AC99
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1), .IN1(~na267_1), .IN2(na272_1), .IN3(~na271_1), .IN4(na250_1), .IN5(1'b0), .IN6(na251_1), .IN7(na216_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y81     80'h00_0018_00_0000_0666_A9CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(1'b0), .IN2(na3475_1), .IN3(1'b0), .IN4(na269_1), .IN5(~na268_1), .IN6(na3475_2), .IN7(na256_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y81     80'h00_0018_00_0040_0AD1_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_1 ( .OUT(na268_1), .IN1(1'b1), .IN2(na239_1), .IN3(1'b1), .IN4(~na218_1), .IN5(~na3478_2), .IN6(1'b0), .IN7(na240_2),
                     .IN8(na248_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x82y82     80'h00_0018_00_0040_0AD3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_1 ( .OUT(na269_1), .IN1(~na244_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na245_1), .IN5(~na246_1), .IN6(1'b1), .IN7(na3485_1),
                     .IN8(na4186_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x82y83     80'h00_0018_00_0040_0AB2_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_1 ( .OUT(na271_1), .IN1(1'b1), .IN2(~na4188_2), .IN3(1'b1), .IN4(na4185_2), .IN5(na246_1), .IN6(~na3467_1), .IN7(1'b0),
                     .IN8(na248_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x83y84     80'h00_0018_00_0040_0CC7_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1), .IN1(na3487_2), .IN2(na3477_2), .IN3(~na240_2), .IN4(1'b1), .IN5(~na244_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na218_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x92y83     80'h00_0018_00_0000_0666_A65C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1), .IN1(1'b0), .IN2(na255_1), .IN3(~na254_1), .IN4(1'b0), .IN5(~na252_1), .IN6(~na259_1), .IN7(na260_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x137y72     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a274_1 ( .OUT(na274_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3489_1), .IN6(~na275_1), .IN7(1'b0), .IN8(~na25_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y74     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a275_1 ( .OUT(na275_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3490_2), .IN6(~na1134_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x123y82     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a276_4 ( .OUT(na276_2), .IN1(~na21_1), .IN2(~na2052_1), .IN3(~na2020_1), .IN4(na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x118y78     80'h40_E818_00_0000_0666_5A90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na273_1), .IN4(na265_1), .IN5(na215_1), .IN6(1'b0), .IN7(~na278_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a277_5 ( .OUT(na277_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na277_1) );
// C_XOR////      x90y67     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na267_1), .IN6(1'b0), .IN7(1'b0), .IN8(na249_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x146y65     80'h40_E800_00_0000_0788_EF35
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a279_1 ( .OUT(na279_1_i), .IN1(~na283_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na280_1), .IN5(1'b1), .IN6(1'b1), .IN7(na3494_1),
                     .IN8(na25_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a279_2 ( .OUT(na279_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na279_1_i) );
// C_MX4b////      x140y78     80'h00_0018_00_0040_0AA0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_1 ( .OUT(na280_1), .IN1(~na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1451_2), .IN5(1'b0), .IN6(na1989_2), .IN7(1'b0), .IN8(na277_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x133y75     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3496_1), .IN6(~na1135_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x141y71     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1451_2), .IN5(1'b0), .IN6(~na285_1), .IN7(1'b0), .IN8(~na3497_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y80     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2920_2), .IN6(na4192_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x129y84     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_1 ( .OUT(na285_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_1), .IN6(~na2053_2), .IN7(~na2021_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x116y61     80'h40_E818_00_0000_0666_9A5A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1), .IN1(na215_2), .IN2(1'b0), .IN3(~na278_1), .IN4(1'b0), .IN5(na215_1), .IN6(1'b0), .IN7(na273_1),
                     .IN8(~na249_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a287_5 ( .OUT(na287_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na287_1) );
// C_MX4b////      x84y87     80'h00_0018_00_0040_0A74_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a290_1 ( .OUT(na290_1), .IN1(~na244_1), .IN2(1'b1), .IN3(1'b1), .IN4(na245_1), .IN5(na3501_1), .IN6(na4190_2), .IN7(~na225_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y86     80'h00_0018_00_0040_0ABD_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a291_1 ( .OUT(na291_1), .IN1(1'b1), .IN2(~na4179_2), .IN3(1'b1), .IN4(na4185_2), .IN5(~na4187_2), .IN6(na3502_1), .IN7(1'b1),
                     .IN8(~na4106_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x129y66     80'h00_0060_00_0000_0C08_FF3B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a292_4 ( .OUT(na292_2), .IN1(na3504_2), .IN2(~na293_1), .IN3(1'b0), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y68     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a293_1 ( .OUT(na293_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1136_1), .IN8(~na3505_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x124y69     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a294_4 ( .OUT(na294_2), .IN1(~na21_1), .IN2(~na2054_1), .IN3(~na2022_1), .IN4(na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x100y65     80'h40_E818_00_0000_0666_AC9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_1 ( .OUT(na295_1), .IN1(na215_2), .IN2(1'b0), .IN3(na278_1), .IN4(~na249_2), .IN5(1'b0), .IN6(na296_1), .IN7(na273_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a295_5 ( .OUT(na295_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na295_1) );
// C_XOR////      x81y72     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a296_1 ( .OUT(na296_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na267_1), .IN6(na272_1), .IN7(na271_1), .IN8(na249_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x129y66     80'h00_0018_00_0000_0C88_3DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a297_1 ( .OUT(na297_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na298_1), .IN6(na3509_2), .IN7(1'b0), .IN8(~na25_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y67     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a298_1 ( .OUT(na298_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3510_2), .IN6(~na1137_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x119y72     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a299_4 ( .OUT(na299_2), .IN1(~na21_1), .IN2(~na2055_2), .IN3(~na2023_2), .IN4(na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x121y61     80'h40_E818_00_0000_0666_500C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a300_1 ( .OUT(na300_1), .IN1(1'b0), .IN2(na303_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na301_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a300_5 ( .OUT(na300_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na300_1) );
// C_///XOR/      x90y61     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a301_4 ( .OUT(na301_2), .IN1(na215_2), .IN2(~na296_1), .IN3(na216_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x81y68     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a303_4 ( .OUT(na303_2), .IN1(na268_1), .IN2(1'b0), .IN3(1'b0), .IN4(na269_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x134y69     80'h00_0018_00_0000_0888_F737
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a304_1 ( .OUT(na304_1), .IN1(~na26_1), .IN2(~na1147_2), .IN3(1'b0), .IN4(~na306_1), .IN5(~na26_2), .IN6(~na2415_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y72     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a306_1 ( .OUT(na306_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na300_2), .IN6(na2923_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y67     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_1 ( .OUT(na307_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3515_1), .IN6(~na1138_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x112y70     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a308_1 ( .OUT(na308_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_1), .IN6(~na2056_1), .IN7(~na2024_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x121y60     80'h40_E818_00_0000_0666_A0C0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na310_1), .IN5(1'b0), .IN6(1'b0), .IN7(na301_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a309_5 ( .OUT(na309_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na309_1) );
// C_XOR////      x90y64     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a310_1 ( .OUT(na310_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na278_1), .IN8(~na265_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y65     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2924_2), .IN6(na309_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x126y61     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_1 ( .OUT(na312_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3519_2), .IN6(~na313_1), .IN7(1'b0), .IN8(~na25_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y64     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a313_1 ( .OUT(na313_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1139_1), .IN8(~na3520_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x128y62     80'h00_0060_00_0000_0C08_FFD7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a314_4 ( .OUT(na314_2), .IN1(~na21_1), .IN2(~na2057_2), .IN3(~na2025_2), .IN4(na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x111y61     80'h40_E818_00_0000_0666_A9CA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a315_1 ( .OUT(na315_1), .IN1(na215_2), .IN2(1'b0), .IN3(1'b0), .IN4(na265_1), .IN5(na215_1), .IN6(~na296_1), .IN7(na216_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a315_5 ( .OUT(na315_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na315_1) );
// C_ORAND*/D///      x136y59     80'h40_E800_00_0000_0788_EF55
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a316_1 ( .OUT(na316_1_i), .IN1(~na320_1), .IN2(1'b0), .IN3(~na317_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3524_2),
                     .IN8(na25_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a316_2 ( .OUT(na316_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na316_1_i) );
// C_MX4b////      x124y59     80'h00_0018_00_0040_0A50_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a317_1 ( .OUT(na317_1), .IN1(na21_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(na315_1), .IN6(1'b0), .IN7(na1994_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y61     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3526_2), .IN8(~na1140_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y59     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_1 ( .OUT(na320_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na3527_2), .IN7(1'b0), .IN8(~na322_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y68     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na315_2), .IN6(na2925_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y62     80'h00_0018_00_0000_0C88_D7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_1), .IN6(~na2058_1), .IN7(~na2026_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x137y63     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na325_1), .IN6(1'b0), .IN7(~na330_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a324_2 ( .OUT(na324_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na324_1_i) );
// C_AND////      x133y73     80'h00_0018_00_0000_0888_54F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(~na3531_2), .IN2(~na328_1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3531_1), .IN6(na329_1), .IN7(~na327_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y79     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2942_2), .IN6(na1077_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y78     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1109_1),
                     .IN8(na2379_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y80     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na861_1), .IN8(~na2402_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x116y79     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a330_1 ( .OUT(na330_1), .IN1(~na21_1), .IN2(~na2043_2), .IN3(~na2107_2), .IN4(na25_1), .IN5(na21_2), .IN6(~na1979_2), .IN7(~na2011_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x148y65     80'h40_E800_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a333_1 ( .OUT(na333_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1451_2), .IN5(~na339_1), .IN6(1'b0), .IN7(~na334_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a333_2 ( .OUT(na333_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na333_1_i) );
// C_AND////      x130y83     80'h00_0018_00_0000_0888_231F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a334_1 ( .OUT(na334_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na337_1), .IN4(~na3536_2), .IN5(1'b1), .IN6(~na336_1), .IN7(na338_1),
                     .IN8(~na3536_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y80     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a336_1 ( .OUT(na336_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na1078_1), .IN6(na2943_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y81     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a337_1 ( .OUT(na337_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1110_1),
                     .IN8(na2380_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y79     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a338_1 ( .OUT(na338_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na870_1), .IN8(~na2403_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x127y85     80'h00_0018_00_0000_0888_D7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a339_1 ( .OUT(na339_1), .IN1(na21_2), .IN2(~na1980_1), .IN3(~na2108_1), .IN4(na25_1), .IN5(~na21_1), .IN6(~na2044_1), .IN7(~na2012_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x147y65     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a342_1 ( .OUT(na342_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na343_1), .IN6(1'b0), .IN7(~na350_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a342_2 ( .OUT(na342_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na342_1_i) );
// C_AND////      x141y77     80'h00_0018_00_0000_0888_1552
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(na3543_2), .IN2(~na3541_1), .IN3(~na3544_1), .IN4(1'b1), .IN5(~na346_1), .IN6(1'b1), .IN7(~na3544_2),
                     .IN8(~na345_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y84     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a345_1 ( .OUT(na345_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na1079_1), .IN6(na2944_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y79     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a346_1 ( .OUT(na346_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1111_1),
                     .IN8(na2381_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x144y77     80'h00_0078_00_0000_0C88_3C33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1333_2), .IN7(1'b1), .IN8(~na25_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a349_4 ( .OUT(na349_2), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x132y85     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a350_1 ( .OUT(na350_1), .IN1(~na21_1), .IN2(~na2045_1), .IN3(~na2109_2), .IN4(na25_1), .IN5(na21_2), .IN6(~na1981_2), .IN7(~na2013_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x142y59     80'h40_E800_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1451_2), .IN5(~na359_1), .IN6(1'b0), .IN7(~na354_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a353_2 ( .OUT(na353_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na353_1_i) );
// C_AND////      x142y69     80'h00_0018_00_0000_0888_1332
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(na3550_2), .IN2(~na3548_2), .IN3(1'b1), .IN4(~na3551_1), .IN5(1'b1), .IN6(~na357_1), .IN7(~na356_1),
                     .IN8(~na3551_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x130y77     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na1080_1), .IN6(na2945_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y72     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na1112_1), .IN6(na2382_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x121y73     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1), .IN1(~na21_1), .IN2(~na2046_1), .IN3(~na2110_1), .IN4(na25_1), .IN5(na21_2), .IN6(~na1982_1), .IN7(~na2014_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x134y61     80'h40_E800_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_1 ( .OUT(na362_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na363_1), .IN7(1'b0), .IN8(~na368_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a362_2 ( .OUT(na362_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na362_1_i) );
// C_AND////      x127y70     80'h00_0018_00_0000_0888_4555
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1), .IN1(~na366_1), .IN2(1'b1), .IN3(~na4381_2), .IN4(1'b1), .IN5(~na3555_1), .IN6(1'b1), .IN7(~na365_1),
                     .IN8(na367_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y73     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a365_1 ( .OUT(na365_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2946_2), .IN8(na1081_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y75     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na2383_2), .IN6(na1113_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y74     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_1 ( .OUT(na367_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na886_1), .IN8(~na2406_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x116y72     80'h00_0018_00_0000_0888_D7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_1 ( .OUT(na368_1), .IN1(na21_2), .IN2(~na1983_2), .IN3(~na2111_2), .IN4(na25_1), .IN5(~na21_1), .IN6(~na2047_2), .IN7(~na2015_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x114y68     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a371_1 ( .OUT(na371_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na3560_1), .IN6(1'b0), .IN7(~na374_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a371_2 ( .OUT(na371_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na371_1_i) );
// C_ORAND////      x104y71     80'h00_0018_00_0000_0888_7BDB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_1 ( .OUT(na374_1), .IN1(na4174_2), .IN2(~na2112_1), .IN3(~na2016_1), .IN4(na25_2), .IN5(na21_2), .IN6(~na1984_2), .IN7(~na2048_1),
                     .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y73     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1082_1), .IN8(na2947_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y71     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_1 ( .OUT(na379_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1114_1),
                     .IN8(na2384_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x132y60     80'h40_E800_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a380_1 ( .OUT(na380_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1451_2), .IN5(1'b0), .IN6(~na386_1), .IN7(1'b0), .IN8(~na381_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a380_2 ( .OUT(na380_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na380_1_i) );
// C_AND////      x140y66     80'h00_0018_00_0000_0888_1545
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1), .IN1(~na3572_1), .IN2(1'b1), .IN3(~na3569_1), .IN4(na3571_2), .IN5(~na3572_2), .IN6(1'b1), .IN7(~na383_1),
                     .IN8(~na384_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y71     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a383_1 ( .OUT(na383_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2948_2), .IN8(na1083_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y70     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a384_1 ( .OUT(na384_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1115_1),
                     .IN8(na2385_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x121y64     80'h00_0018_00_0000_0888_D7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(na21_2), .IN2(~na1985_2), .IN3(~na2113_2), .IN4(na25_1), .IN5(~na21_1), .IN6(~na2049_2), .IN7(~na2017_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x135y60     80'h40_E800_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a389_1 ( .OUT(na389_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1451_2), .IN5(~na3576_1), .IN6(1'b0), .IN7(~na390_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a389_2 ( .OUT(na389_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na389_1_i) );
// C_AND////      x130y63     80'h00_0018_00_0000_0888_3132
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a390_1 ( .OUT(na390_1), .IN1(na3579_1), .IN2(~na3580_1), .IN3(1'b1), .IN4(~na3577_1), .IN5(~na392_1), .IN6(~na3580_2), .IN7(1'b1),
                     .IN8(~na393_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y69     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a392_1 ( .OUT(na392_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2949_1), .IN6(na1084_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y68     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1116_1),
                     .IN8(na2386_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x146y66     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a397_1 ( .OUT(na397_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na398_1), .IN6(1'b0), .IN7(~na3585_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a397_2 ( .OUT(na397_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na397_1_i) );
// C_AND////      x153y93     80'h00_0018_00_0000_0888_5134
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a398_1 ( .OUT(na398_1), .IN1(~na3589_1), .IN2(na3588_2), .IN3(1'b1), .IN4(~na3586_1), .IN5(~na3589_2), .IN6(~na401_1), .IN7(~na400_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y93     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a400_1 ( .OUT(na400_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1085_1), .IN8(na2371_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y92     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a401_1 ( .OUT(na401_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1117_1),
                     .IN8(na2426_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x150y72     80'h40_E800_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a405_1 ( .OUT(na405_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na406_1), .IN7(1'b0), .IN8(~na411_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a405_2 ( .OUT(na405_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na405_1_i) );
// C_AND////      x149y94     80'h00_0018_00_0000_0888_2533
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a406_1 ( .OUT(na406_1), .IN1(1'b1), .IN2(~na409_1), .IN3(1'b1), .IN4(~na3594_2), .IN5(~na408_1), .IN6(1'b1), .IN7(na410_1),
                     .IN8(~na3594_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y91     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na1086_1), .IN6(na2372_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y94     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a409_1 ( .OUT(na409_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na2427_1), .IN6(na1118_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y93     80'h00_0018_00_0040_0A3F_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a410_1 ( .OUT(na410_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(~na940_2), .IN6(~na948_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x128y88     80'h00_0018_00_0000_0888_D7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(na21_2), .IN2(~na1972_1), .IN3(~na2068_1), .IN4(na25_1), .IN5(~na21_1), .IN6(~na2036_1), .IN7(~na2004_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x151y66     80'h40_E800_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a414_1 ( .OUT(na414_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na415_1), .IN7(1'b0), .IN8(~na420_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a414_2 ( .OUT(na414_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na414_1_i) );
// C_AND////      x151y92     80'h00_0018_00_0000_0888_1554
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1), .IN1(~na3599_1), .IN2(na3601_2), .IN3(~na3602_2), .IN4(1'b1), .IN5(~na417_1), .IN6(1'b1), .IN7(~na3602_1),
                     .IN8(~na418_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y89     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2373_2), .IN8(na1087_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y88     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a418_1 ( .OUT(na418_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1119_1),
                     .IN8(na2428_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x130y86     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a420_1 ( .OUT(na420_1), .IN1(~na21_1), .IN2(~na2037_2), .IN3(~na2069_2), .IN4(na25_1), .IN5(na21_2), .IN6(~na1973_2), .IN7(~na2005_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x145y64     80'h40_E800_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na3606_1), .IN7(1'b0), .IN8(~na426_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a423_2 ( .OUT(na423_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na423_1_i) );
// C_ORAND////      x122y76     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a426_1 ( .OUT(na426_1), .IN1(~na21_1), .IN2(~na2038_1), .IN3(~na2070_1), .IN4(na25_1), .IN5(na21_2), .IN6(~na1974_1), .IN7(~na2006_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y90     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_1 ( .OUT(na430_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2374_1), .IN8(na1088_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y87     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1), .IN1(1'b1), .IN2(na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2429_2),
                     .IN8(na1120_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x139y64     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a432_1 ( .OUT(na432_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na3614_1), .IN6(1'b0), .IN7(~na433_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a432_2 ( .OUT(na432_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na432_1_i) );
// C_ORAND////      x116y73     80'h00_0018_00_0000_0888_7BDD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a433_1 ( .OUT(na433_1), .IN1(~na2071_2), .IN2(na4175_2), .IN3(~na2007_2), .IN4(na25_2), .IN5(na21_2), .IN6(~na1975_2), .IN7(~na2039_2),
                     .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y89     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na962_2), .IN8(~na964_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y83     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_1 ( .OUT(na439_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1089_1), .IN8(na2375_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y86     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_1 ( .OUT(na440_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1121_1),
                     .IN8(na2430_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x119y63     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a441_1 ( .OUT(na441_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na442_1), .IN6(1'b0), .IN7(~na3621_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a441_2 ( .OUT(na441_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na441_1_i) );
// C_AND////      x151y89     80'h00_0018_00_0000_0888_3154
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1), .IN1(~na3625_1), .IN2(na3624_1), .IN3(~na3622_2), .IN4(1'b1), .IN5(~na3625_2), .IN6(~na444_1), .IN7(1'b1),
                     .IN8(~na445_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y96     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a444_1 ( .OUT(na444_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1090_1), .IN8(na2376_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x146y86     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a445_1 ( .OUT(na445_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na2431_1), .IN6(na1122_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x136y62     80'h40_E800_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_1 ( .OUT(na449_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na450_1), .IN7(1'b0), .IN8(~na455_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a449_2 ( .OUT(na449_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na449_1_i) );
// C_AND////      x151y82     80'h00_0018_00_0000_0888_1323
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a450_1 ( .OUT(na450_1), .IN1(1'b1), .IN2(~na3633_2), .IN3(na3632_1), .IN4(~na3630_2), .IN5(1'b1), .IN6(~na3633_1), .IN7(~na452_1),
                     .IN8(~na453_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y79     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na1091_1), .IN6(na2377_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x140y82     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a453_1 ( .OUT(na453_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na2432_2), .IN6(na1123_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x114y66     80'h00_0018_00_0000_0888_D7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1), .IN1(na21_2), .IN2(~na1977_2), .IN3(~na2073_2), .IN4(na25_1), .IN5(~na21_1), .IN6(~na2041_2), .IN7(~na2009_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x134y65     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a458_1 ( .OUT(na458_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na3637_1), .IN6(1'b0), .IN7(~na461_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a458_2 ( .OUT(na458_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na458_1_i) );
// C_ORAND////      x122y65     80'h00_0018_00_0000_0888_7BDB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_1 ( .OUT(na461_1), .IN1(na4174_2), .IN2(~na2074_1), .IN3(~na2010_1), .IN4(na25_2), .IN5(na21_2), .IN6(~na1978_1), .IN7(~na2042_1),
                     .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x143y77     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na1092_1), .IN6(na2378_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y76     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na2433_1), .IN6(na1124_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x146y67     80'h40_E800_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1451_2), .IN5(1'b0), .IN6(~na473_1), .IN7(1'b0), .IN8(~na468_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a467_2 ( .OUT(na467_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na467_1_i) );
// C_AND////      x142y84     80'h00_0018_00_0000_0888_2F15
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a468_1 ( .OUT(na468_1), .IN1(~na471_1), .IN2(1'b1), .IN3(~na4382_2), .IN4(~na3646_1), .IN5(1'b1), .IN6(1'b1), .IN7(na472_1),
                     .IN8(~na470_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x132y90     80'h00_0018_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na1093_1), .IN6(na2418_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x137y87     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_1 ( .OUT(na471_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1125_1),
                     .IN8(na972_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y89     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a472_1 ( .OUT(na472_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1017_1),
                     .IN8(~na2926_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x117y80     80'h00_0018_00_0000_0888_D7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a473_1 ( .OUT(na473_1), .IN1(na21_2), .IN2(~na3198_1), .IN3(~na2059_2), .IN4(na25_1), .IN5(~na21_1), .IN6(~na2027_2), .IN7(~na1995_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x149y67     80'h40_E800_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_1 ( .OUT(na476_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1451_2), .IN5(1'b0), .IN6(~na477_1), .IN7(1'b0), .IN8(~na3651_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a476_2 ( .OUT(na476_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na476_1_i) );
// C_ORAND////      x139y96     80'h00_0018_00_0000_0888_7BDD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1), .IN1(~na2060_1), .IN2(na4175_2), .IN3(~na1996_1), .IN4(na25_2), .IN5(na21_2), .IN6(~na3199_2), .IN7(~na2028_1),
                     .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x139y80     80'h00_0060_00_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a481_4 ( .OUT(na481_2), .IN1(~na21_1), .IN2(na3657_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x134y88     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a483_1 ( .OUT(na483_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2419_1), .IN8(na1094_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y83     80'h00_0018_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_1 ( .OUT(na484_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na1126_1), .IN6(na1018_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x150y68     80'h40_E800_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a485_1 ( .OUT(na485_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1451_2), .IN5(~na491_1), .IN6(1'b0), .IN7(~na486_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a485_2 ( .OUT(na485_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na485_1_i) );
// C_AND////      x152y89     80'h00_0018_00_0000_0888_311A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1), .IN1(na3661_1), .IN2(1'b1), .IN3(~na4384_2), .IN4(~na3662_2), .IN5(~na3659_2), .IN6(~na488_1), .IN7(1'b1),
                     .IN8(~na489_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y90     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a488_1 ( .OUT(na488_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1095_1), .IN8(na2420_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y90     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_1 ( .OUT(na489_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na4309_2), .IN6(na1127_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x129y85     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1), .IN1(~na21_1), .IN2(~na2029_2), .IN3(~na2061_2), .IN4(na25_1), .IN5(na21_2), .IN6(~na3200_1), .IN7(~na1997_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x142y64     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a494_1 ( .OUT(na494_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na495_1), .IN6(1'b0), .IN7(~na500_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a494_2 ( .OUT(na494_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na494_1_i) );
// C_AND////      x147y81     80'h00_0018_00_0000_0888_1352
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1), .IN1(na3668_2), .IN2(~na3669_1), .IN3(~na3666_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na3669_2), .IN7(~na497_1),
                     .IN8(~na498_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y87     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_1 ( .OUT(na497_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2421_1), .IN6(na1096_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y86     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a498_1 ( .OUT(na498_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na4311_2), .IN6(na1128_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y73     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a500_1 ( .OUT(na500_1), .IN1(~na21_1), .IN2(~na2030_1), .IN3(~na2062_1), .IN4(na25_1), .IN5(na21_2), .IN6(~na3201_2), .IN7(~na1998_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x137y61     80'h40_E800_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(~na504_1), .IN6(1'b0), .IN7(~na509_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a503_2 ( .OUT(na503_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na503_1_i) );
// C_AND////      x149y81     80'h00_0018_00_0000_0888_4353
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a504_1 ( .OUT(na504_1), .IN1(1'b1), .IN2(~na3673_1), .IN3(~na507_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3673_2), .IN7(~na506_1),
                     .IN8(na508_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x138y85     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a506_1 ( .OUT(na506_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2422_2), .IN6(na1097_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y85     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a507_1 ( .OUT(na507_1), .IN1(1'b1), .IN2(na1333_2), .IN3(na4173_2), .IN4(1'b1), .IN5(na1041_2), .IN6(na1129_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x134y80     80'h00_0060_00_0000_0C0E_FF5A
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a508_4 ( .OUT(na508_2), .IN1(na3675_1), .IN2(1'b0), .IN3(~na4171_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x116y75     80'h00_0018_00_0000_0888_D7DB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a509_1 ( .OUT(na509_1), .IN1(na21_2), .IN2(~na3202_1), .IN3(~na2063_2), .IN4(na25_1), .IN5(~na21_1), .IN6(~na2031_2), .IN7(~na1999_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x123y62     80'h40_E800_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a512_1 ( .OUT(na512_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na3679_1), .IN7(1'b0), .IN8(~na515_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a512_2 ( .OUT(na512_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na512_1_i) );
// C_ORAND////      x106y72     80'h00_0018_00_0000_0888_7BDD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a515_1 ( .OUT(na515_1), .IN1(~na2064_1), .IN2(na4175_2), .IN3(~na2000_1), .IN4(na25_2), .IN5(na21_2), .IN6(~na3203_2), .IN7(~na2032_1),
                     .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y83     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a519_1 ( .OUT(na519_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2423_1), .IN6(na1098_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y84     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a520_1 ( .OUT(na520_1), .IN1(1'b1), .IN2(na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1045_2),
                     .IN8(na1130_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x131y60     80'h40_E800_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a521_1 ( .OUT(na521_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1451_2), .IN5(~na527_1), .IN6(1'b0), .IN7(~na522_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a521_2 ( .OUT(na521_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na521_1_i) );
// C_AND////      x142y71     80'h00_0018_00_0000_0888_5123
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a522_1 ( .OUT(na522_1), .IN1(1'b1), .IN2(~na3691_2), .IN3(na3690_1), .IN4(~na3688_2), .IN5(~na524_1), .IN6(~na3691_1), .IN7(~na525_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y79     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a524_1 ( .OUT(na524_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2424_2), .IN8(na1099_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y77     80'h00_0018_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1131_1),
                     .IN8(na1049_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x113y65     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a527_1 ( .OUT(na527_1), .IN1(~na21_1), .IN2(~na2033_2), .IN3(~na2065_2), .IN4(na25_1), .IN5(na21_2), .IN6(~na3204_1), .IN7(~na2001_2),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x133y59     80'h40_E800_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a530_1 ( .OUT(na530_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(~na531_1), .IN7(1'b0), .IN8(~na536_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a530_2 ( .OUT(na530_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na530_1_i) );
// C_AND////      x145y72     80'h00_0018_00_0000_0888_341F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a531_1 ( .OUT(na531_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na534_1), .IN4(~na3695_1), .IN5(~na533_1), .IN6(na535_1), .IN7(1'b1),
                     .IN8(~na3695_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x131y77     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(na25_2), .IN5(na2425_1), .IN6(na1100_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y75     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a534_1 ( .OUT(na534_1), .IN1(1'b1), .IN2(na1333_2), .IN3(~na4173_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1051_2),
                     .IN8(na1132_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x133y76     80'h00_0018_00_0040_0A3F_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a535_1 ( .OUT(na535_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(na25_1), .IN5(~na1052_1), .IN6(~na2933_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y64     80'h00_0018_00_0000_0888_DBD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a536_1 ( .OUT(na536_1), .IN1(~na21_1), .IN2(~na2034_1), .IN3(~na2066_1), .IN4(na25_1), .IN5(na21_2), .IN6(~na3205_2), .IN7(~na2002_1),
                     .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*/D///      x145y59     80'h40_EC00_00_0000_0388_2FFF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a539_1 ( .OUT(na539_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na540_1), .IN8(~na544_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a539_2 ( .OUT(na539_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na539_1_i) );
// C_MX4b////      x126y59     80'h00_0018_00_0040_0A3B_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a540_1 ( .OUT(na540_1), .IN1(na539_1), .IN2(1'b1), .IN3(1'b1), .IN4(na549_1), .IN5(~na542_2), .IN6(~na541_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x125y60     80'h00_0018_00_0040_0CF3_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a541_1 ( .OUT(na541_1), .IN1(~na1331_1), .IN2(~na3700_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1859_1), .IN7(1'b1),
                     .IN8(na1332_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y75     80'h00_0060_00_0000_0C08_FFC8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a542_4 ( .OUT(na542_2), .IN1(na6_1), .IN2(na5_1), .IN3(1'b1), .IN4(na543_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x84y76     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a543_4 ( .OUT(na543_2), .IN1(~na3_1), .IN2(~na5_2), .IN3(~na2_1), .IN4(~na4165_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x146y60     80'h00_0018_00_0000_0C88_42FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a544_1 ( .OUT(na544_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na539_1), .IN6(~na545_2), .IN7(~na3701_1), .IN8(na549_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x149y66     80'h00_0060_00_0000_0C08_FF18
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a545_4 ( .OUT(na545_2), .IN1(na546_2), .IN2(na12_1), .IN3(~na4166_2), .IN4(~na9_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x153y65     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a546_4 ( .OUT(na546_2), .IN1(~na10_1), .IN2(~na12_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y60     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a547_1 ( .OUT(na547_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3235_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1386_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND*/D      x149y59     80'h40_E800_80_0000_0C07_FFCA
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a548_4 ( .OUT(na548_2_i), .IN1(na539_1), .IN2(1'b1), .IN3(1'b1), .IN4(na549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a548_5 ( .OUT(na548_2), .CLK(1'b0), .EN(na549_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na548_2_i) );
// C_MX2b/D///      x146y62     80'h40_EC00_00_0040_0A54_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a549_1 ( .OUT(na549_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na549_1), .IN5(na3702_1), .IN6(1'b0), .IN7(~na550_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a549_2 ( .OUT(na549_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na549_1_i) );
// C_AND////      x150y61     80'h00_0018_00_0000_0C88_58FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a550_1 ( .OUT(na550_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na539_1), .IN6(na545_2), .IN7(~na3701_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x95y90     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a551_1 ( .OUT(na551_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2203_2), .IN6(na1582_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a551_2 ( .OUT(na551_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na551_1_i) );
// C_///OR/      x113y75     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a552_4 ( .OUT(na552_2), .IN1(~na3294_2), .IN2(~na1859_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x111y83     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a553_1 ( .OUT(na553_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1583_1), .IN6(na2204_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a553_2 ( .OUT(na553_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na553_1_i) );
// C_MX2b/D///      x111y92     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a554_1 ( .OUT(na554_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2205_2), .IN8(na1584_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a554_2 ( .OUT(na554_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na554_1_i) );
// C_MX2b/D///      x107y67     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a555_1 ( .OUT(na555_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1585_1), .IN6(na2206_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a555_2 ( .OUT(na555_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na555_1_i) );
// C_MX2b/D///      x97y75     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a556_1 ( .OUT(na556_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1586_1), .IN6(na2207_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a556_2 ( .OUT(na556_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na556_1_i) );
// C_MX2b/D///      x81y74     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a557_1 ( .OUT(na557_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1587_2), .IN6(na2208_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a557_2 ( .OUT(na557_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na557_1_i) );
// C_MX2b/D///      x93y63     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a558_1 ( .OUT(na558_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1588_2), .IN6(na2209_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a558_2 ( .OUT(na558_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na558_1_i) );
// C_MX2b/D///      x98y63     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a559_1 ( .OUT(na559_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1589_1), .IN8(na2210_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a559_2 ( .OUT(na559_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na559_1_i) );
// C_MX2b/D///      x95y91     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a560_1 ( .OUT(na560_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2211_2), .IN6(na1590_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a560_2 ( .OUT(na560_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na560_1_i) );
// C_MX2b/D///      x107y89     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a561_1 ( .OUT(na561_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1591_1), .IN6(na2212_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a561_2 ( .OUT(na561_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na561_1_i) );
// C_MX2b/D///      x103y96     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a562_1 ( .OUT(na562_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2213_2), .IN6(na1592_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a562_2 ( .OUT(na562_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na562_1_i) );
// C_MX2b/D///      x101y75     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a563_1 ( .OUT(na563_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1593_1), .IN6(na2214_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a563_2 ( .OUT(na563_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na563_1_i) );
// C_MX2b/D///      x91y79     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a564_1 ( .OUT(na564_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2215_2), .IN8(na1594_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a564_2 ( .OUT(na564_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na564_1_i) );
// C_MX2b/D///      x83y73     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a565_1 ( .OUT(na565_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1595_2), .IN6(na2216_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a565_2 ( .OUT(na565_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na565_1_i) );
// C_MX2b/D///      x88y67     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a566_1 ( .OUT(na566_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1596_1), .IN8(na2217_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a566_2 ( .OUT(na566_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na566_1_i) );
// C_MX2b/D///      x92y66     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2218_1), .IN6(na1597_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a567_2 ( .OUT(na567_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na567_1_i) );
// C_MX2b/D///      x121y95     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a568_1 ( .OUT(na568_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2219_2), .IN6(na1598_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a568_2 ( .OUT(na568_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na568_1_i) );
// C_MX2b/D///      x125y97     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_1 ( .OUT(na569_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2220_1), .IN6(na1599_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a569_2 ( .OUT(na569_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na569_1_i) );
// C_MX2b/D///      x123y97     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a570_1 ( .OUT(na570_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1600_1), .IN6(na2221_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a570_2 ( .OUT(na570_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na570_1_i) );
// C_MX2b/D///      x125y91     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a571_1 ( .OUT(na571_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1601_2), .IN8(na2222_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a571_2 ( .OUT(na571_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na571_1_i) );
// C_MX2b/D///      x117y85     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a572_1 ( .OUT(na572_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1602_2), .IN6(na2223_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a572_2 ( .OUT(na572_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na572_1_i) );
// C_MX2b/D///      x107y88     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a573_1 ( .OUT(na573_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2224_1), .IN6(na1603_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a573_2 ( .OUT(na573_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na573_1_i) );
// C_MX2b/D///      x106y66     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a574_1 ( .OUT(na574_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1604_2), .IN8(na2225_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a574_2 ( .OUT(na574_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na574_1_i) );
// C_MX2b/D///      x115y69     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a575_1 ( .OUT(na575_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2226_1), .IN6(na1605_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a575_2 ( .OUT(na575_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na575_1_i) );
// C_MX2b/D///      x105y93     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a576_1 ( .OUT(na576_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1606_2), .IN6(na2171_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a576_2 ( .OUT(na576_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na576_1_i) );
// C_MX2b/D///      x112y95     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_1 ( .OUT(na577_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1607_1), .IN8(na2172_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a577_2 ( .OUT(na577_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na577_1_i) );
// C_MX2b/D///      x116y95     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a578_1 ( .OUT(na578_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2173_2), .IN8(na1608_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a578_2 ( .OUT(na578_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na578_1_i) );
// C_MX2b/D///      x105y87     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_1 ( .OUT(na579_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1609_1), .IN6(na2174_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a579_2 ( .OUT(na579_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na579_1_i) );
// C_MX2b/D///      x99y89     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a580_1 ( .OUT(na580_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2175_2), .IN6(na1610_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a580_2 ( .OUT(na580_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na580_1_i) );
// C_MX2b/D///      x94y87     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_1 ( .OUT(na581_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1611_2), .IN6(na2176_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a581_2 ( .OUT(na581_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na581_1_i) );
// C_MX2b/D///      x90y69     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a582_1 ( .OUT(na582_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2177_2), .IN6(na1612_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a582_2 ( .OUT(na582_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na582_1_i) );
// C_MX2b/D///      x92y69     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_1 ( .OUT(na583_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1613_2), .IN6(na2178_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a583_2 ( .OUT(na583_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na583_1_i) );
// C_MX2b/D///      x99y93     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a584_1 ( .OUT(na584_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1734_1), .IN6(na3206_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a584_2 ( .OUT(na584_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na584_1_i) );
// C_MX2b/D///      x111y94     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_1 ( .OUT(na585_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1735_1), .IN6(na3207_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a585_2 ( .OUT(na585_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na585_1_i) );
// C_MX2b/D///      x113y95     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a586_1 ( .OUT(na586_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1736_1), .IN6(na3208_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a586_2 ( .OUT(na586_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na586_1_i) );
// C_MX2b/D///      x101y84     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_1 ( .OUT(na587_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1737_2), .IN6(na3209_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a587_2 ( .OUT(na587_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na587_1_i) );
// C_MX2b/D///      x98y90     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a588_1 ( .OUT(na588_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3210_1), .IN6(na1738_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a588_2 ( .OUT(na588_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na588_1_i) );
// C_MX2b/D///      x89y85     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a589_1 ( .OUT(na589_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1739_1), .IN8(na3211_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a589_2 ( .OUT(na589_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na589_1_i) );
// C_MX2b/D///      x87y68     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a590_1 ( .OUT(na590_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1740_2), .IN6(na3212_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a590_2 ( .OUT(na590_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na590_1_i) );
// C_MX2b/D///      x96y70     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a591_1 ( .OUT(na591_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3213_2), .IN6(na1741_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a591_2 ( .OUT(na591_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na591_1_i) );
// C_MX2b/D///      x97y91     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a592_1 ( .OUT(na592_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3154_2), .IN6(na1710_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a592_2 ( .OUT(na592_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na592_1_i) );
// C_MX2b/D///      x113y86     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a593_1 ( .OUT(na593_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1711_1), .IN6(na3155_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a593_2 ( .OUT(na593_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na593_1_i) );
// C_MX2b/D///      x111y91     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_1 ( .OUT(na594_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1712_1), .IN6(na3156_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a594_2 ( .OUT(na594_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na594_1_i) );
// C_MX2b/D///      x107y70     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a595_1 ( .OUT(na595_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1713_1), .IN8(na3157_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a595_2 ( .OUT(na595_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na595_1_i) );
// C_MX2b/D///      x99y76     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a596_1 ( .OUT(na596_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1714_1), .IN8(na3158_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a596_2 ( .OUT(na596_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na596_1_i) );
// C_MX2b/D///      x83y75     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a597_1 ( .OUT(na597_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1715_1), .IN6(na3159_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a597_2 ( .OUT(na597_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na597_1_i) );
// C_MX2b/D///      x88y65     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a598_1 ( .OUT(na598_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1716_1), .IN6(na3160_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a598_2 ( .OUT(na598_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na598_1_i) );
// C_MX2b/D///      x101y63     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a599_1 ( .OUT(na599_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1717_1), .IN6(na3161_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a599_2 ( .OUT(na599_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na599_1_i) );
// C_MX2b/D///      x99y94     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a600_1 ( .OUT(na600_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1924_2), .IN6(na1718_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a600_2 ( .OUT(na600_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na600_1_i) );
// C_MX2b/D///      x115y92     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a601_1 ( .OUT(na601_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1925_1), .IN6(na1719_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a601_2 ( .OUT(na601_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na601_1_i) );
// C_MX2b/D///      x109y95     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a602_1 ( .OUT(na602_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1926_2), .IN6(na1720_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a602_2 ( .OUT(na602_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na602_1_i) );
// C_MX2b/D///      x110y81     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a603_1 ( .OUT(na603_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1721_1), .IN6(na1927_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a603_2 ( .OUT(na603_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na603_1_i) );
// C_MX2b/D///      x97y76     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a604_1 ( .OUT(na604_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1722_2), .IN6(na1928_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a604_2 ( .OUT(na604_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na604_1_i) );
// C_MX2b/D///      x91y81     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a605_1 ( .OUT(na605_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1723_2), .IN6(na1929_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a605_2 ( .OUT(na605_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na605_1_i) );
// C_MX2b/D///      x91y67     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a606_1 ( .OUT(na606_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1724_2), .IN8(na1930_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a606_2 ( .OUT(na606_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na606_1_i) );
// C_MX2b/D///      x97y68     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a607_1 ( .OUT(na607_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1931_1), .IN8(na1725_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a607_2 ( .OUT(na607_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na607_1_i) );
// C_MX2b/D///      x115y98     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a608_1 ( .OUT(na608_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1726_1), .IN6(na1915_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a608_2 ( .OUT(na608_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na608_1_i) );
// C_MX2b/D///      x125y98     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a609_1 ( .OUT(na609_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1916_2), .IN6(na1727_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a609_2 ( .OUT(na609_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na609_1_i) );
// C_MX2b/D///      x122y98     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a610_1 ( .OUT(na610_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1728_2), .IN8(na1917_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a610_2 ( .OUT(na610_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na610_1_i) );
// C_MX2b/D///      x115y94     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a611_1 ( .OUT(na611_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1918_2), .IN8(na1729_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a611_2 ( .OUT(na611_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na611_1_i) );
// C_MX2b/D///      x111y88     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a612_1 ( .OUT(na612_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1730_1), .IN8(na1919_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a612_2 ( .OUT(na612_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na612_1_i) );
// C_MX2b/D///      x99y83     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a613_1 ( .OUT(na613_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1731_1), .IN8(na1920_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a613_2 ( .OUT(na613_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na613_1_i) );
// C_MX2b/D///      x97y69     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a614_1 ( .OUT(na614_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1921_2), .IN6(na1732_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a614_2 ( .OUT(na614_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na614_1_i) );
// C_MX2b/D///      x110y68     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a615_1 ( .OUT(na615_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1733_2), .IN6(na1922_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a615_2 ( .OUT(na615_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na615_1_i) );
// C_MX2b/D///      x86y78     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a616_1 ( .OUT(na616_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1494_2), .IN8(na2083_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a616_2 ( .OUT(na616_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na616_1_i) );
// C_MX2b/D///      x114y81     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a617_1 ( .OUT(na617_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1495_2), .IN8(na2084_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a617_2 ( .OUT(na617_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na617_1_i) );
// C_MX2b/D///      x115y87     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a618_1 ( .OUT(na618_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1496_1), .IN8(na2085_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a618_2 ( .OUT(na618_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na618_1_i) );
// C_MX2b/D///      x109y62     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a619_1 ( .OUT(na619_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2086_1), .IN8(na1497_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a619_2 ( .OUT(na619_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na619_1_i) );
// C_MX2b/D///      x94y64     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a620_1 ( .OUT(na620_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2087_2), .IN6(na1498_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a620_2 ( .OUT(na620_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na620_1_i) );
// C_MX2b/D///      x85y67     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a621_1 ( .OUT(na621_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2088_1), .IN8(na1499_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a621_2 ( .OUT(na621_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na621_1_i) );
// C_MX2a/D///      x92y61     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a622_1 ( .OUT(na622_1_i), .IN1(na4354_2), .IN2(na2089_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a622_2 ( .OUT(na622_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na622_1_i) );
// C_MX2b/D///      x99y62     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a623_1 ( .OUT(na623_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2090_1), .IN6(na1501_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a623_2 ( .OUT(na623_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na623_1_i) );
// C_MX2a/D///      x88y84     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a624_1 ( .OUT(na624_1_i), .IN1(na2091_2), .IN2(na1502_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a624_2 ( .OUT(na624_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na624_1_i) );
// C_MX2b/D///      x101y89     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a625_1 ( .OUT(na625_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2092_1), .IN8(na1503_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a625_2 ( .OUT(na625_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na625_1_i) );
// C_MX2b/D///      x96y92     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a626_1 ( .OUT(na626_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2093_2), .IN8(na1504_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a626_2 ( .OUT(na626_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na626_1_i) );
// C_MX2b/D///      x101y71     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a627_1 ( .OUT(na627_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2094_1), .IN8(na1505_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a627_2 ( .OUT(na627_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na627_1_i) );
// C_MX2b/D///      x94y73     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a628_1 ( .OUT(na628_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2095_2), .IN6(na1506_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a628_2 ( .OUT(na628_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na628_1_i) );
// C_MX2a/D///      x82y74     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a629_1 ( .OUT(na629_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1507_2), .IN4(na2096_1), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a629_2 ( .OUT(na629_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na629_1_i) );
// C_MX2b/D///      x84y64     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a630_1 ( .OUT(na630_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2097_2), .IN8(na1508_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a630_2 ( .OUT(na630_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na630_1_i) );
// C_MX2a/D///      x87y64     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a631_1 ( .OUT(na631_1_i), .IN1(na1509_2), .IN2(na2098_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a631_2 ( .OUT(na631_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na631_1_i) );
// C_MX2b/D///      x133y99     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a632_1 ( .OUT(na632_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1510_2), .IN8(na1961_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a632_2 ( .OUT(na632_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na632_1_i) );
// C_MX2b/D///      x135y100     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a633_1 ( .OUT(na633_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1511_1), .IN6(na1962_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a633_2 ( .OUT(na633_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na633_1_i) );
// C_MX2b/D///      x127y97     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a634_1 ( .OUT(na634_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1963_2), .IN6(na1512_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a634_2 ( .OUT(na634_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na634_1_i) );
// C_MX2b/D///      x142y94     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1964_1), .IN8(na4355_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a635_2 ( .OUT(na635_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na635_1_i) );
// C_MX2a/D///      x127y84     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a636_1 ( .OUT(na636_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1514_1), .IN4(na1965_2), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a636_2 ( .OUT(na636_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na636_1_i) );
// C_MX2b/D///      x108y82     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a637_1 ( .OUT(na637_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1515_1), .IN6(na1966_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a637_2 ( .OUT(na637_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na637_1_i) );
// C_MX2a/D///      x108y63     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a638_1 ( .OUT(na638_1_i), .IN1(na1967_2), .IN2(na1516_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a638_2 ( .OUT(na638_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na638_1_i) );
// C_MX2b/D///      x124y61     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_1 ( .OUT(na639_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1517_2), .IN8(na1968_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a639_2 ( .OUT(na639_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na639_1_i) );
// C_MX2b/D///      x104y94     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a640_1 ( .OUT(na640_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4353_2), .IN8(na3237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a640_2 ( .OUT(na640_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na640_1_i) );
// C_MX2b/D///      x109y94     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_1 ( .OUT(na641_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1483_2), .IN6(na3238_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a641_2 ( .OUT(na641_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na641_1_i) );
// C_MX2b/D///      x114y96     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a642_1 ( .OUT(na642_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1484_2), .IN6(na3239_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a642_2 ( .OUT(na642_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na642_1_i) );
// C_MX2a/D///      x103y89     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a643_1 ( .OUT(na643_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1486_2), .IN4(na3240_2), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a643_2 ( .OUT(na643_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na643_1_i) );
// C_MX2b/D///      x100y90     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a644_1 ( .OUT(na644_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1488_2), .IN8(na3241_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a644_2 ( .OUT(na644_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na644_1_i) );
// C_MX2a/D///      x84y92     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a645_1 ( .OUT(na645_1_i), .IN1(na1490_2), .IN2(na3242_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a645_2 ( .OUT(na645_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na645_1_i) );
// C_MX2b/D///      x90y76     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a646_1 ( .OUT(na646_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3243_1), .IN8(na1492_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a646_2 ( .OUT(na646_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na646_1_i) );
// C_MX2b/D///      x93y70     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a647_1 ( .OUT(na647_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3244_2), .IN6(na1493_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a647_2 ( .OUT(na647_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na647_1_i) );
// C_MX2b/D///      x93y89     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a648_1 ( .OUT(na648_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2155_2), .IN6(na1518_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a648_2 ( .OUT(na648_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na648_1_i) );
// C_MX2b/D///      x116y82     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a649_1 ( .OUT(na649_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2156_1), .IN6(na1519_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a649_2 ( .OUT(na649_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na649_1_i) );
// C_MX2a/D///      x118y89     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a650_1 ( .OUT(na650_1_i), .IN1(na1520_1), .IN2(na2157_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a650_2 ( .OUT(na650_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na650_1_i) );
// C_MX2b/D///      x113y63     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a651_1 ( .OUT(na651_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2158_1), .IN6(na1521_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a651_2 ( .OUT(na651_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na651_1_i) );
// C_MX2a/D///      x91y65     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a652_1 ( .OUT(na652_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1522_2), .IN4(na2159_2), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a652_2 ( .OUT(na652_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na652_1_i) );
// C_MX2b/D///      x83y67     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a653_1 ( .OUT(na653_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1523_2), .IN6(na2160_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a653_2 ( .OUT(na653_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na653_1_i) );
// C_MX2b/D///      x88y60     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a654_1 ( .OUT(na654_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2161_2), .IN8(na1524_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a654_2 ( .OUT(na654_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na654_1_i) );
// C_MX2b/D///      x100y62     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1525_2), .IN8(na2162_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a655_2 ( .OUT(na655_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na655_1_i) );
// C_MX2b/D///      x92y86     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a656_1 ( .OUT(na656_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2163_2), .IN6(na1526_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a656_2 ( .OUT(na656_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na656_1_i) );
// C_MX2a/D///      x108y92     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a657_1 ( .OUT(na657_1_i), .IN1(na1527_1), .IN2(na2164_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a657_2 ( .OUT(na657_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na657_1_i) );
// C_MX2b/D///      x97y95     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a658_1 ( .OUT(na658_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1528_1), .IN6(na2165_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a658_2 ( .OUT(na658_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na658_1_i) );
// C_MX2a/D///      x97y80     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a659_1 ( .OUT(na659_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1529_2), .IN4(na2166_1), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a659_2 ( .OUT(na659_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na659_1_i) );
// C_MX2b/D///      x89y80     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a660_1 ( .OUT(na660_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2167_1), .IN6(na1530_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a660_2 ( .OUT(na660_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na660_1_i) );
// C_MX2b/D///      x82y76     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a661_1 ( .OUT(na661_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2168_1), .IN6(na1531_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a661_2 ( .OUT(na661_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na661_1_i) );
// C_MX2b/D///      x81y63     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a662_1 ( .OUT(na662_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1532_2), .IN6(na2169_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a662_2 ( .OUT(na662_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na662_1_i) );
// C_MX2b/D///      x88y61     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a663_1 ( .OUT(na663_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2170_1), .IN8(na1533_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a663_2 ( .OUT(na663_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na663_1_i) );
// C_MX2a/D///      x123y96     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a664_1 ( .OUT(na664_1_i), .IN1(na2115_2), .IN2(na1534_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a664_2 ( .OUT(na664_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na664_1_i) );
// C_MX2b/D///      x127y101     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a665_1 ( .OUT(na665_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1535_2), .IN8(na2116_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a665_2 ( .OUT(na665_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na665_1_i) );
// C_MX2a/D///      x122y102     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a666_1 ( .OUT(na666_1_i), .IN1(na1536_1), .IN2(na2117_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a666_2 ( .OUT(na666_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na666_1_i) );
// C_MX2b/D///      x134y93     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a667_1 ( .OUT(na667_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1537_1), .IN6(na2118_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a667_2 ( .OUT(na667_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na667_1_i) );
// C_MX2b/D///      x126y89     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a668_1 ( .OUT(na668_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2119_2), .IN6(na1538_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a668_2 ( .OUT(na668_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na668_1_i) );
// C_MX2b/D///      x109y86     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a669_1 ( .OUT(na669_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1539_2), .IN6(na2120_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a669_2 ( .OUT(na669_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na669_1_i) );
// C_MX2b/D///      x103y61     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a670_1 ( .OUT(na670_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1540_1), .IN6(na2121_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a670_2 ( .OUT(na670_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na670_1_i) );
// C_MX2a/D///      x123y72     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a671_1 ( .OUT(na671_1_i), .IN1(na1541_2), .IN2(na2122_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a671_2 ( .OUT(na671_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na671_1_i) );
// C_MX2b/D///      x110y98     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a672_1 ( .OUT(na672_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2075_2), .IN6(na1542_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a672_2 ( .OUT(na672_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na672_1_i) );
// C_MX2a/D///      x117y100     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a673_1 ( .OUT(na673_1_i), .IN1(na2076_1), .IN2(na1543_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a673_2 ( .OUT(na673_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na673_1_i) );
// C_MX2b/D///      x117y104     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a674_1 ( .OUT(na674_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2077_2), .IN6(na1544_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a674_2 ( .OUT(na674_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na674_1_i) );
// C_MX2b/D///      x105y90     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a675_1 ( .OUT(na675_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2078_1), .IN6(na1545_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a675_2 ( .OUT(na675_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na675_1_i) );
// C_MX2b/D///      x95y94     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a676_1 ( .OUT(na676_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1546_2), .IN6(na2079_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a676_2 ( .OUT(na676_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na676_1_i) );
// C_MX2b/D///      x90y86     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a677_1 ( .OUT(na677_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1547_1), .IN8(na2080_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a677_2 ( .OUT(na677_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na677_1_i) );
// C_MX2a/D///      x85y69     80'h40_E800_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a678_1 ( .OUT(na678_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na2081_2), .IN4(na1548_1), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a678_2 ( .OUT(na678_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na678_1_i) );
// C_MX2b/D///      x89y67     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a679_1 ( .OUT(na679_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2082_1), .IN6(na1549_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a679_2 ( .OUT(na679_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na679_1_i) );
// C_MX2a/D///      x92y88     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a680_1 ( .OUT(na680_1_i), .IN1(na1550_1), .IN2(na2123_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a680_2 ( .OUT(na680_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na680_1_i) );
// C_MX2b/D///      x117y84     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a681_1 ( .OUT(na681_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1551_1), .IN8(na2124_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a681_2 ( .OUT(na681_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na681_1_i) );
// C_MX2b/D///      x119y90     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a682_1 ( .OUT(na682_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2125_2), .IN6(na1552_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a682_2 ( .OUT(na682_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na682_1_i) );
// C_MX2b/D///      x112y64     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a683_1 ( .OUT(na683_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1553_1), .IN8(na2126_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a683_2 ( .OUT(na683_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na683_1_i) );
// C_MX2b/D///      x101y70     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a684_1 ( .OUT(na684_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1554_1), .IN6(na2127_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a684_2 ( .OUT(na684_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na684_1_i) );
// C_MX2a/D///      x86y69     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1_i), .IN1(na2128_1), .IN2(na1555_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a685_2 ( .OUT(na685_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na685_1_i) );
// C_MX2b/D///      x91y62     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a686_1 ( .OUT(na686_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1556_1), .IN8(na2129_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a686_2 ( .OUT(na686_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na686_1_i) );
// C_MX2a/D///      x100y59     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a687_1 ( .OUT(na687_1_i), .IN1(na1557_1), .IN2(na2130_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a687_2 ( .OUT(na687_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na687_1_i) );
// C_MX2b/D///      x92y89     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a688_1 ( .OUT(na688_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1558_2), .IN6(na2131_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a688_2 ( .OUT(na688_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na688_1_i) );
// C_MX2b/D///      x110y91     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a689_1 ( .OUT(na689_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2132_1), .IN6(na1559_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a689_2 ( .OUT(na689_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na689_1_i) );
// C_MX2b/D///      x102y95     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a690_1 ( .OUT(na690_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2133_2), .IN6(na1560_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a690_2 ( .OUT(na690_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na690_1_i) );
// C_MX2b/D///      x94y78     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a691_1 ( .OUT(na691_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2134_1), .IN6(na1561_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a691_2 ( .OUT(na691_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na691_1_i) );
// C_MX2a/D///      x88y77     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a692_1 ( .OUT(na692_1_i), .IN1(na1562_2), .IN2(na2135_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a692_2 ( .OUT(na692_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na692_1_i) );
// C_MX2b/D///      x85y74     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a693_1 ( .OUT(na693_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1563_2), .IN6(na2136_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a693_2 ( .OUT(na693_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na693_1_i) );
// C_MX2a/D///      x87y66     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a694_1 ( .OUT(na694_1_i), .IN1(na1564_1), .IN2(na2137_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a694_2 ( .OUT(na694_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na694_1_i) );
// C_MX2b/D///      x91y64     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1565_2), .IN6(na2138_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a695_2 ( .OUT(na695_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na695_1_i) );
// C_MX2b/D///      x126y95     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a696_1 ( .OUT(na696_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1566_2), .IN8(na2139_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a696_2 ( .OUT(na696_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na696_1_i) );
// C_MX2b/D///      x126y100     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a697_1 ( .OUT(na697_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1567_1), .IN6(na2140_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a697_2 ( .OUT(na697_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na697_1_i) );
// C_MX2b/D///      x130y101     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a698_1 ( .OUT(na698_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1568_1), .IN8(na2141_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a698_2 ( .OUT(na698_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na698_1_i) );
// C_MX2a/D///      x122y92     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a699_1 ( .OUT(na699_1_i), .IN1(na2142_1), .IN2(na1569_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a699_2 ( .OUT(na699_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na699_1_i) );
// C_MX2b/D///      x118y83     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a700_1 ( .OUT(na700_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1570_2), .IN6(na2143_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a700_2 ( .OUT(na700_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na700_1_i) );
// C_MX2a/D///      x102y89     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a701_1 ( .OUT(na701_1_i), .IN1(na2144_1), .IN2(na1571_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a701_2 ( .OUT(na701_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na701_1_i) );
// C_MX2b/D///      x107y62     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2145_2), .IN6(na1572_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a702_2 ( .OUT(na702_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na702_1_i) );
// C_MX2b/D///      x122y67     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1573_1), .IN6(na2146_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a703_2 ( .OUT(na703_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na703_1_i) );
// C_MX2b/D///      x108y95     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a704_1 ( .OUT(na704_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1574_1), .IN6(na2147_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a704_2 ( .OUT(na704_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na704_1_i) );
// C_MX2b/D///      x118y98     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a705_1 ( .OUT(na705_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1575_2), .IN8(na2148_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a705_2 ( .OUT(na705_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na705_1_i) );
// C_MX2a/D///      x120y100     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a706_1 ( .OUT(na706_1_i), .IN1(na1576_1), .IN2(na2149_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a706_2 ( .OUT(na706_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na706_1_i) );
// C_MX2b/D///      x106y90     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1577_2), .IN6(na2150_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a707_2 ( .OUT(na707_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na707_1_i) );
// C_MX2a/D///      x92y92     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a708_1 ( .OUT(na708_1_i), .IN1(na1578_1), .IN2(na2151_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a708_2 ( .OUT(na708_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na708_1_i) );
// C_MX2b/D///      x89y86     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1579_2), .IN6(na2152_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a709_2 ( .OUT(na709_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na709_1_i) );
// C_MX2b/D///      x89y68     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a710_1 ( .OUT(na710_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2153_2), .IN6(na1580_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a710_2 ( .OUT(na710_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na710_1_i) );
// C_MX2b/D///      x90y66     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1581_2), .IN6(na2154_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a711_2 ( .OUT(na711_1), .CLK(1'b0), .EN(na1473_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na711_1_i) );
// C_MX2b/D///      x95y86     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a712_1 ( .OUT(na712_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1614_2), .IN8(na2227_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a712_2 ( .OUT(na712_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na712_1_i) );
// C_MX2a/D///      x123y90     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a713_1 ( .OUT(na713_1_i), .IN1(na1615_1), .IN2(na2228_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a713_2 ( .OUT(na713_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na713_1_i) );
// C_MX2b/D///      x115y90     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a714_1 ( .OUT(na714_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2229_2), .IN6(na1616_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a714_2 ( .OUT(na714_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na714_1_i) );
// C_MX2a/D///      x114y62     80'h40_E800_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a715_1 ( .OUT(na715_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na2230_1), .IN4(na1617_1), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a715_2 ( .OUT(na715_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na715_1_i) );
// C_MX2b/D///      x94y66     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a716_1 ( .OUT(na716_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1618_2), .IN6(na2231_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a716_2 ( .OUT(na716_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na716_1_i) );
// C_MX2b/D///      x85y70     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a717_1 ( .OUT(na717_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1619_2), .IN8(na2232_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a717_2 ( .OUT(na717_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na717_1_i) );
// C_MX2b/D///      x90y62     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a718_1 ( .OUT(na718_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2233_2), .IN6(na4357_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a718_2 ( .OUT(na718_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na718_1_i) );
// C_MX2b/D///      x102y60     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1621_2), .IN6(na2234_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a719_2 ( .OUT(na719_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na719_1_i) );
// C_MX2a/D///      x93y91     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a720_1 ( .OUT(na720_1_i), .IN1(na1622_2), .IN2(na2179_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a720_2 ( .OUT(na720_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na720_1_i) );
// C_MX2b/D///      x107y93     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2180_1), .IN6(na1623_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a721_2 ( .OUT(na721_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na721_1_i) );
// C_MX2a/D///      x101y96     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a722_1 ( .OUT(na722_1_i), .IN1(na2181_2), .IN2(na4358_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a722_2 ( .OUT(na722_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na722_1_i) );
// C_MX2b/D///      x106y76     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1625_1), .IN6(na2182_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a723_2 ( .OUT(na723_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na723_1_i) );
// C_MX2b/D///      x96y77     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a724_1 ( .OUT(na724_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2183_2), .IN6(na1626_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a724_2 ( .OUT(na724_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na724_1_i) );
// C_MX2b/D///      x85y80     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a725_1 ( .OUT(na725_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2184_1), .IN6(na1627_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a725_2 ( .OUT(na725_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na725_1_i) );
// C_MX2b/D///      x87y65     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a726_1 ( .OUT(na726_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1628_2), .IN8(na2185_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a726_2 ( .OUT(na726_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na726_1_i) );
// C_MX2a/D///      x89y66     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1_i), .IN1(na1629_2), .IN2(na2186_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a727_2 ( .OUT(na727_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na727_1_i) );
// C_MX2b/D///      x128y95     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a728_1 ( .OUT(na728_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2187_2), .IN8(na1630_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a728_2 ( .OUT(na728_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na728_1_i) );
// C_MX2a/D///      x129y102     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a729_1 ( .OUT(na729_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1631_2), .IN4(na2188_1), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a729_2 ( .OUT(na729_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na729_1_i) );
// C_MX2b/D///      x128y98     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a730_1 ( .OUT(na730_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1632_2), .IN6(na2189_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a730_2 ( .OUT(na730_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na730_1_i) );
// C_MX2b/D///      x129y92     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1633_2), .IN6(na2190_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a731_2 ( .OUT(na731_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na731_1_i) );
// C_MX2b/D///      x129y94     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a732_1 ( .OUT(na732_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1634_2), .IN6(na2191_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a732_2 ( .OUT(na732_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na732_1_i) );
// C_MX2b/D///      x115y82     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a733_1 ( .OUT(na733_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1635_2), .IN6(na2192_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a733_2 ( .OUT(na733_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na733_1_i) );
// C_MX2a/D///      x104y64     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a734_1 ( .OUT(na734_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1636_2), .IN4(na2193_2), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a734_2 ( .OUT(na734_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na734_1_i) );
// C_MX2b/D///      x122y72     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a735_1 ( .OUT(na735_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2194_1), .IN8(na1637_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a735_2 ( .OUT(na735_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na735_1_i) );
// C_MX2a/D///      x108y96     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a736_1 ( .OUT(na736_1_i), .IN1(na2195_2), .IN2(na4359_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a736_2 ( .OUT(na736_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na736_1_i) );
// C_MX2b/D///      x111y96     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1639_2), .IN6(na2196_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a737_2 ( .OUT(na737_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na737_1_i) );
// C_MX2b/D///      x125y100     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a738_1 ( .OUT(na738_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2197_2), .IN6(na1640_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a738_2 ( .OUT(na738_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na738_1_i) );
// C_MX2b/D///      x103y91     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1641_2), .IN6(na2198_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a739_2 ( .OUT(na739_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na739_1_i) );
// C_MX2b/D///      x101y92     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a740_1 ( .OUT(na740_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1642_2), .IN8(na2199_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a740_2 ( .OUT(na740_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na740_1_i) );
// C_MX2a/D///      x89y94     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a741_1 ( .OUT(na741_1_i), .IN1(na2200_1), .IN2(na1643_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a741_2 ( .OUT(na741_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na741_1_i) );
// C_MX2b/D///      x101y69     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a742_1 ( .OUT(na742_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1644_2), .IN8(na2201_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a742_2 ( .OUT(na742_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na742_1_i) );
// C_MX2a/D///      x105y70     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a743_1 ( .OUT(na743_1_i), .IN1(na1645_1), .IN2(na2202_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a743_2 ( .OUT(na743_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na743_1_i) );
// C_MX2b/D///      x93y90     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a744_1 ( .OUT(na744_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1646_1), .IN6(na2251_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a744_2 ( .OUT(na744_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na744_1_i) );
// C_MX2b/D///      x124y89     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a745_1 ( .OUT(na745_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1647_2), .IN6(na2252_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a745_2 ( .OUT(na745_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na745_1_i) );
// C_MX2b/D///      x117y93     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a746_1 ( .OUT(na746_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2253_2), .IN6(na1648_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a746_2 ( .OUT(na746_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na746_1_i) );
// C_MX2b/D///      x115y63     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a747_1 ( .OUT(na747_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1649_2), .IN6(na2254_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a747_2 ( .OUT(na747_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na747_1_i) );
// C_MX2a/D///      x95y68     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a748_1 ( .OUT(na748_1_i), .IN1(na2255_2), .IN2(na1650_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a748_2 ( .OUT(na748_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na748_1_i) );
// C_MX2b/D///      x84y72     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a749_1 ( .OUT(na749_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1651_1), .IN6(na2256_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a749_2 ( .OUT(na749_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na749_1_i) );
// C_MX2a/D///      x89y59     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a750_1 ( .OUT(na750_1_i), .IN1(na1652_2), .IN2(na2257_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a750_2 ( .OUT(na750_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na750_1_i) );
// C_MX2b/D///      x104y61     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a751_1 ( .OUT(na751_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1653_2), .IN6(na2258_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a751_2 ( .OUT(na751_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na751_1_i) );
// C_MX2b/D///      x88y87     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a752_1 ( .OUT(na752_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1654_2), .IN6(na2259_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a752_2 ( .OUT(na752_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na752_1_i) );
// C_MX2b/D///      x108y93     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_1 ( .OUT(na753_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1655_1), .IN6(na2260_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a753_2 ( .OUT(na753_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na753_1_i) );
// C_MX2b/D///      x100y95     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a754_1 ( .OUT(na754_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2261_2), .IN6(na1656_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a754_2 ( .OUT(na754_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na754_1_i) );
// C_MX2a/D///      x97y81     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a755_1 ( .OUT(na755_1_i), .IN1(na2262_1), .IN2(na1657_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a755_2 ( .OUT(na755_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na755_1_i) );
// C_MX2b/D///      x95y83     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a756_1 ( .OUT(na756_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1658_2), .IN6(na2263_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a756_2 ( .OUT(na756_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na756_1_i) );
// C_MX2a/D///      x84y79     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a757_1 ( .OUT(na757_1_i), .IN1(na2264_1), .IN2(na1659_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a757_2 ( .OUT(na757_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na757_1_i) );
// C_MX2b/D///      x85y64     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a758_1 ( .OUT(na758_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1660_1), .IN6(na2265_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a758_2 ( .OUT(na758_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na758_1_i) );
// C_MX2b/D///      x86y62     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_1 ( .OUT(na759_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1661_1), .IN6(na2266_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a759_2 ( .OUT(na759_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na759_1_i) );
// C_MX2b/D///      x125y99     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a760_1 ( .OUT(na760_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1662_1), .IN8(na2267_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a760_2 ( .OUT(na760_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na760_1_i) );
// C_MX2b/D///      x124y102     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a761_1 ( .OUT(na761_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2268_1), .IN6(na1663_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a761_2 ( .OUT(na761_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na761_1_i) );
// C_MX2a/D///      x129y100     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a762_1 ( .OUT(na762_1_i), .IN1(na1664_2), .IN2(na2269_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a762_2 ( .OUT(na762_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na762_1_i) );
// C_MX2b/D///      x120y96     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a763_1 ( .OUT(na763_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1665_1), .IN8(na2270_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a763_2 ( .OUT(na763_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na763_1_i) );
// C_MX2a/D///      x126y92     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a764_1 ( .OUT(na764_1_i), .IN1(na2271_2), .IN2(na1666_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a764_2 ( .OUT(na764_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na764_1_i) );
// C_MX2b/D///      x103y85     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1667_2), .IN8(na2272_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a765_2 ( .OUT(na765_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na765_1_i) );
// C_MX2b/D///      x97y62     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a766_1 ( .OUT(na766_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1668_1), .IN6(na2273_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a766_2 ( .OUT(na766_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na766_1_i) );
// C_MX2b/D///      x125y73     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a767_1 ( .OUT(na767_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2274_1), .IN6(na1669_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a767_2 ( .OUT(na767_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na767_1_i) );
// C_MX2b/D///      x112y97     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a768_1 ( .OUT(na768_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2275_2), .IN6(na1670_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a768_2 ( .OUT(na768_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na768_1_i) );
// C_MX2a/D///      x118y99     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a769_1 ( .OUT(na769_1_i), .IN1(na1671_2), .IN2(na2276_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a769_2 ( .OUT(na769_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na769_1_i) );
// C_MX2b/D///      x120y101     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a770_1 ( .OUT(na770_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2277_2), .IN6(na1672_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a770_2 ( .OUT(na770_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na770_1_i) );
// C_MX2a/D///      x100y92     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a771_1 ( .OUT(na771_1_i), .IN1(na1673_1), .IN2(na2278_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a771_2 ( .OUT(na771_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na771_1_i) );
// C_MX2b/D///      x95y93     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a772_1 ( .OUT(na772_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2279_2), .IN6(na1674_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a772_2 ( .OUT(na772_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na772_1_i) );
// C_MX2b/D///      x87y87     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a773_1 ( .OUT(na773_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2280_1), .IN6(na1675_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a773_2 ( .OUT(na773_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na773_1_i) );
// C_MX2b/D///      x93y76     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a774_1 ( .OUT(na774_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1676_2), .IN6(na2281_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a774_2 ( .OUT(na774_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na774_1_i) );
// C_MX2b/D///      x91y72     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1677_2), .IN6(na2282_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a775_2 ( .OUT(na775_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na775_1_i) );
// C_MX2a/D///      x96y90     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a776_1 ( .OUT(na776_1_i), .IN1(na3165_2), .IN2(na1678_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a776_2 ( .OUT(na776_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na776_1_i) );
// C_MX2b/D///      x120y84     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1679_1), .IN6(na3166_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a777_2 ( .OUT(na777_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na777_1_i) );
// C_MX2a/D///      x118y93     80'h40_E800_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a778_1 ( .OUT(na778_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3167_2), .IN4(na1680_2), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a778_2 ( .OUT(na778_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na778_1_i) );
// C_MX2b/D///      x111y66     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1681_1), .IN6(na3168_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a779_2 ( .OUT(na779_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na779_1_i) );
// C_MX2b/D///      x98y69     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a780_1 ( .OUT(na780_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1682_2), .IN6(na3169_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a780_2 ( .OUT(na780_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na780_1_i) );
// C_MX2b/D///      x85y72     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3170_1), .IN6(na1683_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a781_2 ( .OUT(na781_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na781_1_i) );
// C_MX2b/D///      x89y62     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a782_1 ( .OUT(na782_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3171_2), .IN8(na1684_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a782_2 ( .OUT(na782_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na782_1_i) );
// C_MX2a/D///      x103y62     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1_i), .IN1(na1685_2), .IN2(na3172_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a783_2 ( .OUT(na783_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na783_1_i) );
// C_MX2b/D///      x94y88     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a784_1 ( .OUT(na784_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2283_2), .IN6(na1686_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a784_2 ( .OUT(na784_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na784_1_i) );
// C_MX2a/D///      x106y92     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_1 ( .OUT(na785_1_i), .IN1(na1687_1), .IN2(na2284_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a785_2 ( .OUT(na785_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na785_1_i) );
// C_MX2b/D///      x105y96     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a786_1 ( .OUT(na786_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1688_1), .IN8(na2285_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a786_2 ( .OUT(na786_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na786_1_i) );
// C_MX2b/D///      x100y80     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1689_2), .IN6(na2286_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a787_2 ( .OUT(na787_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na787_1_i) );
// C_MX2b/D///      x96y81     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a788_1 ( .OUT(na788_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2287_2), .IN6(na1690_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a788_2 ( .OUT(na788_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na788_1_i) );
// C_MX2b/D///      x86y80     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1691_2), .IN8(na2288_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a789_2 ( .OUT(na789_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na789_1_i) );
// C_MX2a/D///      x86y64     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a790_1 ( .OUT(na790_1_i), .IN1(na2289_1), .IN2(na1692_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a790_2 ( .OUT(na790_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na790_1_i) );
// C_MX2b/D///      x90y63     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_1 ( .OUT(na791_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1693_2), .IN6(na2290_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a791_2 ( .OUT(na791_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na791_1_i) );
// C_MX2a/D///      x117y96     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a792_1 ( .OUT(na792_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1694_1), .IN4(na2235_2), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a792_2 ( .OUT(na792_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na792_1_i) );
// C_MX2b/D///      x126y101     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a793_1 ( .OUT(na793_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1695_2), .IN6(na2236_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a793_2 ( .OUT(na793_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na793_1_i) );
// C_MX2b/D///      x130y99     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a794_1 ( .OUT(na794_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2237_2), .IN6(na1696_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a794_2 ( .OUT(na794_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na794_1_i) );
// C_MX2b/D///      x132y89     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a795_1 ( .OUT(na795_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2238_1), .IN8(na1697_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a795_2 ( .OUT(na795_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na795_1_i) );
// C_MX2b/D///      x120y89     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_1 ( .OUT(na796_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2239_2), .IN6(na1698_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a796_2 ( .OUT(na796_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na796_1_i) );
// C_MX2a/D///      x106y88     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1_i), .IN1(na1699_1), .IN2(na2240_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a797_2 ( .OUT(na797_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na797_1_i) );
// C_MX2b/D///      x102y62     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a798_1 ( .OUT(na798_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2241_2), .IN6(na1700_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a798_2 ( .OUT(na798_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na798_1_i) );
// C_MX2a/D///      x118y65     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a799_1 ( .OUT(na799_1_i), .IN1(na2242_1), .IN2(na1701_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a799_2 ( .OUT(na799_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na799_1_i) );
// C_MX2b/D///      x109y96     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a800_1 ( .OUT(na800_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1702_1), .IN6(na2243_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a800_2 ( .OUT(na800_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na800_1_i) );
// C_MX2b/D///      x115y96     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a801_1 ( .OUT(na801_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2244_1), .IN8(na1703_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a801_2 ( .OUT(na801_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na801_1_i) );
// C_MX2b/D///      x118y102     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a802_1 ( .OUT(na802_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2245_2), .IN8(na1704_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a802_2 ( .OUT(na802_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na802_1_i) );
// C_MX2b/D///      x102y87     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a803_1 ( .OUT(na803_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1705_2), .IN8(na2246_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a803_2 ( .OUT(na803_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na803_1_i) );
// C_MX2a/D///      x99y90     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a804_1 ( .OUT(na804_1_i), .IN1(na2247_2), .IN2(na1706_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a804_2 ( .OUT(na804_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na804_1_i) );
// C_MX2b/D///      x90y87     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a805_1 ( .OUT(na805_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1707_2), .IN6(na2248_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a805_2 ( .OUT(na805_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na805_1_i) );
// C_MX2a/D///      x90y68     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a806_1 ( .OUT(na806_1_i), .IN1(na1708_1), .IN2(na2249_2), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a806_2 ( .OUT(na806_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na806_1_i) );
// C_MX2b/D///      x91y66     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a807_1 ( .OUT(na807_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2250_1), .IN6(na1709_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a807_2 ( .OUT(na807_1), .CLK(1'b0), .EN(na1475_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na807_1_i) );
// C_///AND/D      x106y99     80'h40_E800_80_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a808_4 ( .OUT(na808_2_i), .IN1(1'b1), .IN2(~na4240_2), .IN3(na809_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a808_5 ( .OUT(na808_2), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na808_2_i) );
// C_AND////D      x110y97     80'h40_E818_00_0000_0888_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a809_5 ( .OUT(na809_2), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na809_1) );
// C_///AND/D      x107y101     80'h40_E800_80_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a810_4 ( .OUT(na810_2_i), .IN1(1'b1), .IN2(~na4240_2), .IN3(na808_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a810_5 ( .OUT(na810_2), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na810_2_i) );
// C_AND/D///      x105y97     80'h40_E800_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a811_1 ( .OUT(na811_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na810_2), .IN6(1'b1), .IN7(~na809_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a811_2 ( .OUT(na811_1), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na811_1_i) );
// C_AND/D///      x97y97     80'h40_E800_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a812_1 ( .OUT(na812_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na811_1), .IN6(1'b1), .IN7(~na809_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a812_2 ( .OUT(na812_1), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na812_1_i) );
// C_AND/D///      x90y96     80'h40_E800_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a813_1 ( .OUT(na813_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na812_1), .IN6(1'b1), .IN7(~na809_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a813_2 ( .OUT(na813_1), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na813_1_i) );
// C_///AND/D      x90y96     80'h40_E800_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a814_4 ( .OUT(na814_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na809_1), .IN4(na813_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a814_5 ( .OUT(na814_2), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na814_2_i) );
// C_AND/D///      x88y86     80'h40_E800_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a815_1 ( .OUT(na815_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na809_1), .IN8(na814_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a815_2 ( .OUT(na815_1), .CLK(1'b0), .EN(na1464_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na815_1_i) );
// C_XOR////D      x115y78     80'h40_E818_00_0000_0666_0C0C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a816_1 ( .OUT(na816_1), .IN1(1'b0), .IN2(na855_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na817_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a816_5 ( .OUT(na816_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na816_1) );
// C_XOR////      x85y82     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na818_2), .IN6(1'b0), .IN7(1'b0), .IN8(na849_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x85y81     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a818_4 ( .OUT(na818_2), .IN1(1'b0), .IN2(1'b0), .IN3(na819_1), .IN4(na843_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y85     80'h00_0018_00_0040_0AD0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a819_1 ( .OUT(na819_1), .IN1(1'b1), .IN2(na820_1), .IN3(~na3705_2), .IN4(1'b1), .IN5(na3723_2), .IN6(1'b0), .IN7(na3705_1),
                     .IN8(na839_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y92     80'h00_0018_00_0040_0AF5_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a820_1 ( .OUT(na820_1), .IN1(~na1842_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4252_2), .IN5(~na3706_1), .IN6(na4385_2), .IN7(~na1844_1),
                     .IN8(na836_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x86y102     80'h00_0078_00_0000_0C66_A9CA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a821_1 ( .OUT(na821_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1168_1), .IN6(na822_2), .IN7(na824_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a821_4 ( .OUT(na821_2), .IN1(na1170_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1172_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x91y102     80'h00_0060_00_0000_0C06_FF56
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a822_4 ( .OUT(na822_2), .IN1(na1178_1), .IN2(na1180_1), .IN3(~na1176_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x88y101     80'h00_0078_00_0000_0C66_905C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a824_1 ( .OUT(na824_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1176_1), .IN8(~na1172_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a824_4 ( .OUT(na824_2), .IN1(1'b0), .IN2(na1180_1), .IN3(~na1176_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x85y101     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a825_1 ( .OUT(na825_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1170_1), .IN6(1'b0), .IN7(na1182_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x90y100     80'h00_0018_00_0040_0A62_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a826_1 ( .OUT(na826_1), .IN1(na1178_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1172_1), .IN5(1'b0), .IN6(~na4323_2), .IN7(na1182_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x85y100     80'h00_0078_00_0000_0C66_9969
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1178_1), .IN6(na1174_1), .IN7(~na1182_1),
                     .IN8(na1172_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a827_4 ( .OUT(na827_2), .IN1(na1170_1), .IN2(~na1180_1), .IN3(na1176_1), .IN4(na4324_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x81y102     80'h00_0018_00_0000_0666_5DDE
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a829_1 ( .OUT(na829_1), .IN1(~na825_1), .IN2(~na822_2), .IN3(na4249_2), .IN4(~na821_1), .IN5(na4244_2), .IN6(~na827_2), .IN7(na832_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y101     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a832_1 ( .OUT(na832_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4386_2), .IN5(na3711_1), .IN6(1'b0), .IN7(na1176_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x84y102     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a834_1 ( .OUT(na834_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na827_2), .IN7(~na824_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x80y102     80'h00_0018_00_0000_0666_C3DA
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a836_1 ( .OUT(na836_1), .IN1(~na4246_2), .IN2(1'b1), .IN3(na4243_2), .IN4(~na4386_2), .IN5(1'b1), .IN6(na838_1), .IN7(1'b1),
                     .IN8(~na3715_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y102     80'h00_0018_00_0040_0A75_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a838_1 ( .OUT(na838_1), .IN1(na1178_1), .IN2(1'b1), .IN3(~na824_2), .IN4(1'b1), .IN5(~na825_1), .IN6(na3716_2), .IN7(~na824_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y90     80'h00_0018_00_0040_0AF2_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_1 ( .OUT(na839_1), .IN1(1'b1), .IN2(na829_1), .IN3(1'b1), .IN4(na836_1), .IN5(na1842_1), .IN6(~na4362_2), .IN7(na1844_1),
                     .IN8(na3717_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x96y99     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a842_4 ( .OUT(na842_2), .IN1(1'b0), .IN2(na1174_1), .IN3(1'b0), .IN4(na1172_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y88     80'h00_0018_00_0040_0A7E_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a843_1 ( .OUT(na843_1), .IN1(1'b1), .IN2(~na844_1), .IN3(1'b1), .IN4(na845_1), .IN5(na3718_2), .IN6(~na846_2), .IN7(~na848_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y98     80'h00_0018_00_0040_0AF8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a844_1 ( .OUT(na844_1), .IN1(na1842_1), .IN2(1'b1), .IN3(~na1844_1), .IN4(1'b1), .IN5(na4253_2), .IN6(na829_1), .IN7(na3719_1),
                     .IN8(~na836_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y94     80'h00_0018_00_0040_0AF5_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a845_1 ( .OUT(na845_1), .IN1(1'b1), .IN2(na829_1), .IN3(na1844_1), .IN4(1'b1), .IN5(~na1842_1), .IN6(na3720_2), .IN7(~na4254_2),
                     .IN8(na836_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x81y100     80'h00_0060_00_0000_0C06_FF3A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a846_4 ( .OUT(na846_2), .IN1(na1168_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na3728_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y97     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a848_1 ( .OUT(na848_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1170_1), .IN6(na827_2), .IN7(1'b0), .IN8(na1172_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y96     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a849_1 ( .OUT(na849_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na852_1), .IN6(na851_1), .IN7(na850_1), .IN8(na853_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x88y97     80'h00_0018_00_0040_0A7A_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a850_1 ( .OUT(na850_1), .IN1(1'b1), .IN2(na820_1), .IN3(1'b1), .IN4(na4386_2), .IN5(na3721_1), .IN6(~na844_1), .IN7(na4245_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y98     80'h00_0018_00_0040_0ABD_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a851_1 ( .OUT(na851_1), .IN1(1'b1), .IN2(~na827_2), .IN3(1'b1), .IN4(na845_1), .IN5(~na4248_2), .IN6(na3722_2), .IN7(1'b1),
                     .IN8(~na839_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y99     80'h00_0018_00_0040_0AB2_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a852_1 ( .OUT(na852_1), .IN1(1'b1), .IN2(na827_1), .IN3(na4251_2), .IN4(1'b1), .IN5(na3723_1), .IN6(~na820_1), .IN7(1'b0),
                     .IN8(na839_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x86y100     80'h00_0018_00_0040_0ADB_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_1 ( .OUT(na853_1), .IN1(1'b1), .IN2(~na844_1), .IN3(1'b1), .IN4(~na845_1), .IN5(~na854_1), .IN6(1'b1), .IN7(na3724_1),
                     .IN8(~na4255_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y101     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a854_1 ( .OUT(na854_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na822_2), .IN7(1'b0), .IN8(na4386_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x83y96     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a855_4 ( .OUT(na855_2), .IN1(na857_1), .IN2(~na860_1), .IN3(na859_1), .IN4(na858_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x89y97     80'h00_0018_00_0000_0C66_E7FF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_1 ( .OUT(na857_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4256_2), .IN6(na827_1), .IN7(~na4251_2), .IN8(~na845_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x90y98     80'h00_0018_00_0040_0C5B_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a858_1 ( .OUT(na858_1), .IN1(~na854_1), .IN2(na822_2), .IN3(1'b1), .IN4(na4386_2), .IN5(1'b1), .IN6(~na820_1), .IN7(1'b1),
                     .IN8(~na839_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x88y99     80'h00_0018_00_0040_0A7E_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a859_1 ( .OUT(na859_1), .IN1(1'b1), .IN2(na820_1), .IN3(1'b1), .IN4(na3728_2), .IN5(na4388_2), .IN6(~na844_1), .IN7(~na4321_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x79y100     80'h00_0018_00_0040_0C7E_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a860_1 ( .OUT(na860_1), .IN1(1'b1), .IN2(~na4387_2), .IN3(~na848_1), .IN4(na3729_2), .IN5(~na4258_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na839_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x128y81     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a861_1 ( .OUT(na861_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4389_2), .IN6(na816_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a861_2 ( .OUT(na861_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na861_1_i) );
// C_XOR////D      x101y88     80'h40_E818_00_0000_0666_5036
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a862_1 ( .OUT(na862_1), .IN1(na818_2), .IN2(na863_2), .IN3(1'b0), .IN4(~na864_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na867_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a862_5 ( .OUT(na862_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na862_1) );
// C_///XOR/      x85y96     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a863_4 ( .OUT(na863_2), .IN1(~na852_1), .IN2(na860_1), .IN3(na859_1), .IN4(~na853_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x82y78     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a864_4 ( .OUT(na864_2), .IN1(~na866_1), .IN2(na851_1), .IN3(na850_1), .IN4(~na4261_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x83y92     80'h00_0018_00_0040_0C17_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a865_1 ( .OUT(na865_1), .IN1(~na3718_2), .IN2(na846_2), .IN3(na848_1), .IN4(1'b0), .IN5(na4258_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na839_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x83y93     80'h00_0018_00_0040_0C5B_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a866_1 ( .OUT(na866_1), .IN1(~na3723_2), .IN2(na3732_2), .IN3(1'b1), .IN4(na3728_2), .IN5(1'b1), .IN6(~na820_1), .IN7(1'b1),
                     .IN8(~na4257_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x88y89     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a867_4 ( .OUT(na867_2), .IN1(na857_1), .IN2(~na4262_2), .IN3(~na868_1), .IN4(na858_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x86y91     80'h00_0018_00_0040_0C2B_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_1 ( .OUT(na868_1), .IN1(na3723_1), .IN2(~na820_1), .IN3(1'b0), .IN4(na839_1), .IN5(na3723_2), .IN6(1'b1), .IN7(~na848_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x84y90     80'h00_0018_00_0040_0AE3_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1), .IN1(1'b1), .IN2(na844_1), .IN3(1'b1), .IN4(~na845_1), .IN5(1'b1), .IN6(~na846_2), .IN7(na3705_2),
                     .IN8(na3734_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x122y83     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_1 ( .OUT(na870_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4390_2), .IN6(na862_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a870_2 ( .OUT(na870_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na870_1_i) );
// C_XOR////D      x121y84     80'h40_E818_00_0000_0666_0A5C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_1 ( .OUT(na871_1), .IN1(1'b0), .IN2(na873_2), .IN3(~na874_1), .IN4(1'b0), .IN5(na872_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a871_5 ( .OUT(na871_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na871_1) );
// C_XOR////      x89y87     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a872_1 ( .OUT(na872_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na857_1), .IN6(na4259_2), .IN7(na4241_2), .IN8(na858_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x83y90     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a873_4 ( .OUT(na873_2), .IN1(na818_2), .IN2(1'b0), .IN3(na867_2), .IN4(na864_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x88y89     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a874_1 ( .OUT(na874_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na875_1), .IN6(na863_2), .IN7(1'b0), .IN8(na849_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x85y81     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_1 ( .OUT(na875_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na868_1), .IN8(na869_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x135y82     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a876_1 ( .OUT(na876_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3736_1), .IN6(na871_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a876_2 ( .OUT(na876_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na876_1_i) );
// C_XOR////D      x123y74     80'h40_E818_00_0000_0666_05C0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_1 ( .OUT(na877_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na878_1), .IN5(~na872_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a877_5 ( .OUT(na877_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na877_1) );
// C_XOR////      x86y86     80'h00_0018_00_0000_0666_6CC9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_1 ( .OUT(na878_1), .IN1(na875_1), .IN2(~na880_1), .IN3(1'b0), .IN4(na869_1), .IN5(1'b0), .IN6(na863_2), .IN7(~na868_1),
                     .IN8(~na881_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y98     80'h00_0018_00_0040_0AE2_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a880_1 ( .OUT(na880_1), .IN1(1'b1), .IN2(na844_1), .IN3(1'b1), .IN4(~na845_1), .IN5(1'b0), .IN6(~na827_2), .IN7(na4260_2),
                     .IN8(na3737_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x84y96     80'h00_0018_00_0040_0C7E_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a881_1 ( .OUT(na881_1), .IN1(1'b1), .IN2(~na827_1), .IN3(~na842_2), .IN4(na3738_1), .IN5(1'b1), .IN6(~na820_1), .IN7(1'b1),
                     .IN8(na839_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x136y74     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a882_1 ( .OUT(na882_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3739_2), .IN6(na877_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a882_2 ( .OUT(na882_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na882_1_i) );
// C_XOR////D      x110y74     80'h40_E818_00_0000_0666_C00C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_1 ( .OUT(na883_1), .IN1(1'b0), .IN2(na884_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na878_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a883_5 ( .OUT(na883_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na883_1) );
// C_///XOR/      x81y86     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a884_4 ( .OUT(na884_2), .IN1(na866_1), .IN2(na865_1), .IN3(na867_2), .IN4(na849_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x124y79     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a886_1 ( .OUT(na886_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3740_1), .IN8(na883_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a886_2 ( .OUT(na886_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na886_1_i) );
// C_XOR////D      x115y72     80'h40_E818_00_0000_0666_AC0A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a887_1 ( .OUT(na887_1), .IN1(na875_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na817_1), .IN7(na888_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a887_5 ( .OUT(na887_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na887_1) );
// C_XOR////      x82y79     80'h00_0018_00_0000_0666_9663
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a888_1 ( .OUT(na888_1), .IN1(1'b0), .IN2(~na880_1), .IN3(na868_1), .IN4(na869_1), .IN5(na866_1), .IN6(na865_1), .IN7(na867_2),
                     .IN8(~na881_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x118y70     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a889_1 ( .OUT(na889_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3741_2), .IN6(na887_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a889_2 ( .OUT(na889_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na889_1_i) );
// C_XOR////D      x124y70     80'h40_E818_00_0000_0666_50C0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a890_1 ( .OUT(na890_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na864_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na888_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a890_5 ( .OUT(na890_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na890_1) );
// C_MX2b/D///      x129y72     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4395_2), .IN8(na890_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a891_2 ( .OUT(na891_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na891_1_i) );
// C_XOR////D      x122y63     80'h40_E818_00_0000_0666_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a892_1 ( .OUT(na892_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na893_2), .IN6(1'b0), .IN7(na888_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a892_5 ( .OUT(na892_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na892_1) );
// C_///XOR/      x85y71     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a893_4 ( .OUT(na893_2), .IN1(na818_2), .IN2(1'b0), .IN3(na4263_2), .IN4(na864_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x124y64     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a894_1 ( .OUT(na894_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na892_1), .IN8(na3743_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a894_2 ( .OUT(na894_1), .CLK(1'b0), .EN(na1453_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na894_1_i) );
// C_XOR////D      x142y98     80'h40_E818_00_0000_0666_A069
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a895_1 ( .OUT(na895_1), .IN1(~na927_1), .IN2(na933_2), .IN3(na896_1), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(na925_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a895_5 ( .OUT(na895_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na895_1) );
// C_XOR////      x146y97     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a896_1 ( .OUT(na896_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na919_1), .IN7(na897_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x154y101     80'h00_0018_00_0040_0ABD_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1), .IN1(~na3744_2), .IN2(1'b1), .IN3(1'b1), .IN4(na898_1), .IN5(~na4325_2), .IN6(na4396_2), .IN7(1'b1),
                     .IN8(~na917_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x156y102     80'h00_0018_00_0040_0AFA_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a898_1 ( .OUT(na898_1), .IN1(1'b1), .IN2(na1847_2), .IN3(na4276_2), .IN4(1'b1), .IN5(na4398_2), .IN6(~na3745_1), .IN7(na3759_2),
                     .IN8(~na911_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y102     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a899_4 ( .OUT(na899_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1198_1), .IN4(~na1186_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y102     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_1 ( .OUT(na900_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1192_1), .IN6(~na1188_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x142y99     80'h00_0078_00_0000_0C66_6669
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a901_1 ( .OUT(na901_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1190_1), .IN6(na1188_1), .IN7(~na1198_1),
                     .IN8(~na1194_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a901_4 ( .OUT(na901_2), .IN1(na1192_1), .IN2(~na1196_1), .IN3(na1198_1), .IN4(na1186_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x144y102     80'h00_0078_00_0000_0C66_56CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a903_1 ( .OUT(na903_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3753_2), .IN6(na900_1), .IN7(~na1184_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a903_4 ( .OUT(na903_2), .IN1(1'b0), .IN2(na1188_1), .IN3(1'b0), .IN4(na1186_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x135y102     80'h00_0018_00_0040_0A64_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a904_1 ( .OUT(na904_1), .IN1(1'b1), .IN2(~na1188_1), .IN3(1'b1), .IN4(na1194_1), .IN5(1'b0), .IN6(na4326_2), .IN7(~na1198_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x143y101     80'h00_0018_00_0000_0666_B5DE
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a906_1 ( .OUT(na906_1), .IN1(~na3753_2), .IN2(~na4269_2), .IN3(na901_1), .IN4(~na903_1), .IN5(na909_1), .IN6(1'b1), .IN7(~na901_2),
                     .IN8(na903_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x139y101     80'h00_0018_00_0000_0C66_B500
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a909_1 ( .OUT(na909_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1192_1), .IN6(1'b1), .IN7(~na3766_2), .IN8(na3750_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y102     80'h00_0018_00_0000_0666_6A06
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a911_1 ( .OUT(na911_1), .IN1(na913_1), .IN2(na914_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3752_1), .IN6(1'b0), .IN7(na1184_1),
                     .IN8(na1194_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x141y101     80'h00_0018_00_0040_0A78_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a913_1 ( .OUT(na913_1), .IN1(na3753_2), .IN2(1'b1), .IN3(na901_2), .IN4(1'b1), .IN5(na3753_1), .IN6(na900_1), .IN7(na1184_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x145y102     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a914_1 ( .OUT(na914_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3766_2), .IN8(na903_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x141y98     80'h00_0060_00_0000_0C08_FF39
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a915_4 ( .OUT(na915_2), .IN1(~na1192_1), .IN2(~na1196_1), .IN3(1'b0), .IN4(na899_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x140y102     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a916_1 ( .OUT(na916_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na901_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1188_1), .IN7(1'b0), .IN8(~na1186_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y102     80'h00_0018_00_0040_0AF4_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a917_1 ( .OUT(na917_1), .IN1(1'b1), .IN2(~na1847_2), .IN3(1'b1), .IN4(~na911_1), .IN5(na906_1), .IN6(na4400_2), .IN7(~na3759_2),
                     .IN8(na3756_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x153y100     80'h00_0018_00_0040_0C7E_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a919_1 ( .OUT(na919_1), .IN1(1'b1), .IN2(~na3768_2), .IN3(~na4280_2), .IN4(na3757_1), .IN5(~na920_1), .IN6(1'b1), .IN7(na921_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x151y101     80'h00_0018_00_0040_0AFA_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_1 ( .OUT(na920_1), .IN1(~na906_1), .IN2(1'b1), .IN3(1'b1), .IN4(na911_1), .IN5(na3758_1), .IN6(~na1847_2), .IN7(na3759_2),
                     .IN8(~na4401_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x156y101     80'h00_0018_00_0040_0AF1_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a921_1 ( .OUT(na921_1), .IN1(~na906_1), .IN2(1'b1), .IN3(na3759_2), .IN4(1'b1), .IN5(~na4363_2), .IN6(na1847_2), .IN7(na3759_1),
                     .IN8(na911_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x142y97     80'h00_0018_00_0000_0C66_7EFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a925_1 ( .OUT(na925_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na920_1), .IN6(~na4274_2), .IN7(na901_1), .IN8(na917_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x144y98     80'h00_0018_00_0040_0CA7_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a926_1 ( .OUT(na926_1), .IN1(na3753_2), .IN2(~na938_1), .IN3(na3766_2), .IN4(1'b1), .IN5(na4268_2), .IN6(1'b1), .IN7(~na921_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y99     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a927_1 ( .OUT(na927_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4402_2), .IN6(na3763_1), .IN7(1'b0), .IN8(na930_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x151y98     80'h00_0078_00_0000_0C66_A59C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a929_1 ( .OUT(na929_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3744_2), .IN6(1'b0), .IN7(na1184_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a929_4 ( .OUT(na929_2), .IN1(1'b0), .IN2(na1188_1), .IN3(na901_2), .IN4(~na1186_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y100     80'h00_0018_00_0040_0A7E_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a930_1 ( .OUT(na930_1), .IN1(na3765_2), .IN2(1'b1), .IN3(1'b1), .IN4(na898_1), .IN5(na3765_1), .IN6(~na3768_2), .IN7(~na921_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y99     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a932_1 ( .OUT(na932_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1190_1), .IN6(na1188_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y100     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a933_4 ( .OUT(na933_2), .IN1(na937_1), .IN2(~na936_1), .IN3(na935_1), .IN4(na4283_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x145y97     80'h00_0018_00_0040_0ADA_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a934_1 ( .OUT(na934_1), .IN1(na4268_2), .IN2(1'b1), .IN3(~na3766_2), .IN4(1'b1), .IN5(na3753_2), .IN6(1'b1), .IN7(na3766_1),
                     .IN8(~na917_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x148y97     80'h00_0018_00_0040_0A7E_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a935_1 ( .OUT(na935_1), .IN1(na920_1), .IN2(1'b1), .IN3(na901_2), .IN4(1'b1), .IN5(na3767_1), .IN6(~na4278_2), .IN7(~na901_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y100     80'h00_0018_00_0040_0A71_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a936_1 ( .OUT(na936_1), .IN1(~na4273_2), .IN2(1'b1), .IN3(na901_2), .IN4(1'b1), .IN5(~na4268_2), .IN6(na3768_1), .IN7(na921_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x147y99     80'h00_0018_00_0040_0ADB_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a937_1 ( .OUT(na937_1), .IN1(na920_1), .IN2(1'b1), .IN3(1'b1), .IN4(na917_1), .IN5(~na932_1), .IN6(1'b1), .IN7(na3769_2),
                     .IN8(~na4284_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y100     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a938_1 ( .OUT(na938_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3753_2), .IN6(1'b0), .IN7(na3766_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x150y94     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a939_1 ( .OUT(na939_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4407_2), .IN8(na895_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a939_2 ( .OUT(na939_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na939_1_i) );
// C_XOR////D      x139y97     80'h40_E818_00_0000_0666_66A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a940_1 ( .OUT(na940_1), .IN1(na943_1), .IN2(~na942_1), .IN3(na925_1), .IN4(1'b0), .IN5(~na937_1), .IN6(~na936_1), .IN7(na896_1),
                     .IN8(na926_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a940_5 ( .OUT(na940_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na940_1) );
// C_XOR////      x145y98     80'h00_0018_00_0000_0666_A9CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a942_1 ( .OUT(na942_1), .IN1(1'b0), .IN2(na3763_2), .IN3(1'b0), .IN4(na930_1), .IN5(~na934_1), .IN6(na3763_1), .IN7(na935_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x151y97     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a943_1 ( .OUT(na943_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na947_1), .IN6(na945_1), .IN7(na944_1), .IN8(~na4286_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x152y97     80'h00_0018_00_0040_0C07_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a944_1 ( .OUT(na944_1), .IN1(na3771_2), .IN2(na929_1), .IN3(na4280_2), .IN4(1'b0), .IN5(na920_1), .IN6(1'b1), .IN7(~na921_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x153y98     80'h00_0018_00_0040_0CA7_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_1 ( .OUT(na945_1), .IN1(na3772_1), .IN2(~na3768_2), .IN3(na4397_2), .IN4(1'b1), .IN5(na4268_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na917_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x155y98     80'h00_0018_00_0040_0C8E_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a946_1 ( .OUT(na946_1), .IN1(1'b0), .IN2(na3768_1), .IN3(na921_1), .IN4(~na898_1), .IN5(1'b1), .IN6(na929_2), .IN7(1'b1),
                     .IN8(na4406_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x153y99     80'h00_0018_00_0040_0A7A_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a947_1 ( .OUT(na947_1), .IN1(na920_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na917_1), .IN5(na3774_2), .IN6(~na929_1), .IN7(na4403_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x139y94     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a948_1 ( .OUT(na948_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4285_2), .IN8(na3775_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a948_2 ( .OUT(na948_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na948_1_i) );
// C_XOR////D      x154y96     80'h40_E818_00_0000_0666_AC50
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a949_1 ( .OUT(na949_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na952_1), .IN4(1'b0), .IN5(1'b0), .IN6(na950_1), .IN7(na951_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a949_5 ( .OUT(na949_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na949_1) );
// C_XOR////      x139y100     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a950_1 ( .OUT(na950_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na927_1), .IN6(na933_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y97     80'h00_0018_00_0000_0666_0969
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a951_1 ( .OUT(na951_1), .IN1(na943_1), .IN2(~na3763_1), .IN3(na935_1), .IN4(na930_1), .IN5(~na934_1), .IN6(na3763_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y99     80'h00_0018_00_0000_0666_666C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a952_1 ( .OUT(na952_1), .IN1(1'b0), .IN2(na933_2), .IN3(~na925_1), .IN4(~na953_2), .IN5(~na937_1), .IN6(~na936_1), .IN7(na896_1),
                     .IN8(na926_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y100     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a953_4 ( .OUT(na953_2), .IN1(~na947_1), .IN2(~na946_1), .IN3(na925_1), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x141y86     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a954_1 ( .OUT(na954_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4409_2), .IN8(na949_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a954_2 ( .OUT(na954_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na954_1_i) );
// C_XOR////D      x143y97     80'h40_E818_00_0000_0666_600A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a955_1 ( .OUT(na955_1), .IN1(na957_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na952_1), .IN8(na956_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a955_5 ( .OUT(na955_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na955_1) );
// C_XOR////      x140y100     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a956_1 ( .OUT(na956_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na927_1), .IN6(~na933_2), .IN7(na925_1), .IN8(na926_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y99     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a957_4 ( .OUT(na957_2), .IN1(na958_2), .IN2(~na933_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x149y97     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a958_4 ( .OUT(na958_2), .IN1(na947_1), .IN2(na946_1), .IN3(~na959_1), .IN4(~na960_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x150y99     80'h00_0018_00_0040_0AE4_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a959_1 ( .OUT(na959_1), .IN1(~na920_1), .IN2(1'b1), .IN3(1'b1), .IN4(na917_1), .IN5(1'b0), .IN6(na938_1), .IN7(~na901_2),
                     .IN8(na3777_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x150y98     80'h00_0018_00_0040_0CE7_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a960_1 ( .OUT(na960_1), .IN1(na3778_2), .IN2(~na4281_2), .IN3(~na901_1), .IN4(1'b1), .IN5(na4268_2), .IN6(1'b1), .IN7(~na921_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x147y93     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a961_1 ( .OUT(na961_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na955_1), .IN6(na3779_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a961_2 ( .OUT(na961_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na961_1_i) );
// C_XOR////D      x154y95     80'h40_E818_00_0000_0666_500A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a962_1 ( .OUT(na962_1), .IN1(na963_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na952_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a962_5 ( .OUT(na962_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na962_1) );
// C_XOR////      x149y95     80'h00_0018_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a963_1 ( .OUT(na963_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na958_2), .IN6(~na945_1), .IN7(~na944_1), .IN8(na953_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x146y90     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a964_1 ( .OUT(na964_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na962_1), .IN8(na4411_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a964_2 ( .OUT(na964_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na964_1_i) );
// C_XOR////D      x153y96     80'h40_E818_00_0000_0666_0AA0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a965_1 ( .OUT(na965_1), .IN1(1'b0), .IN2(1'b0), .IN3(na966_2), .IN4(1'b0), .IN5(na963_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a965_5 ( .OUT(na965_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na965_1) );
// C_///XOR/      x142y101     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a966_4 ( .OUT(na966_2), .IN1(~na947_1), .IN2(~na946_1), .IN3(na4279_2), .IN4(na4282_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x147y86     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a967_1 ( .OUT(na967_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4412_2), .IN6(na965_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a967_2 ( .OUT(na967_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na967_1_i) );
// C_XOR////D      x149y88     80'h40_E818_00_0000_0666_650A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a968_1 ( .OUT(na968_1), .IN1(na958_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na934_1), .IN6(1'b0), .IN7(na935_1), .IN8(na953_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a968_5 ( .OUT(na968_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na968_1) );
// C_MX2b/D///      x147y80     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a969_1 ( .OUT(na969_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4413_2), .IN6(na968_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a969_2 ( .OUT(na969_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na969_1_i) );
// C_XOR////D      x151y81     80'h40_E818_00_0000_0666_A00A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a970_1 ( .OUT(na970_1), .IN1(na963_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na951_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a970_5 ( .OUT(na970_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na970_1) );
// C_MX2b/D///      x143y76     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a971_1 ( .OUT(na971_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na970_1), .IN6(na4414_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a971_2 ( .OUT(na971_1), .CLK(1'b0), .EN(na1456_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na971_1_i) );
// C_XOR////D      x134y94     80'h40_E818_00_0000_0666_030A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a972_1 ( .OUT(na972_1), .IN1(na1014_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na973_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a972_5 ( .OUT(na972_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na972_1) );
// C_XOR////      x115y102     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_1 ( .OUT(na973_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na975_2), .IN6(na999_1), .IN7(na996_1), .IN8(~na4306_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x109y101     80'h00_0060_00_0000_0C06_FFE7
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a975_4 ( .OUT(na975_2), .IN1(na977_1), .IN2(na976_1), .IN3(~na995_1), .IN4(~na4290_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x93y104     80'h00_0018_00_0040_0AF8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a976_1 ( .OUT(na976_1), .IN1(na1852_1), .IN2(1'b1), .IN3(~na989_1), .IN4(1'b1), .IN5(na4418_2), .IN6(na984_1), .IN7(na3786_2),
                     .IN8(~na3800_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x99y99     80'h00_0078_00_0000_0C66_6696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a977_1 ( .OUT(na977_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1210_1), .IN6(~na1214_1), .IN7(na1204_1),
                     .IN8(na1206_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a977_4 ( .OUT(na977_2), .IN1(na1202_1), .IN2(na1214_1), .IN3(~na1212_1), .IN4(na1208_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x98y100     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a978_4 ( .OUT(na978_2), .IN1(~na1202_1), .IN2(na1214_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x97y100     80'h00_0078_00_0000_0C66_9009
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a979_1 ( .OUT(na979_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1204_1), .IN8(na1208_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a979_4 ( .OUT(na979_2), .IN1(~na1210_1), .IN2(na1214_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x96y98     80'h00_0078_00_0000_0C66_C9AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a981_1 ( .OUT(na981_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1200_1), .IN6(na979_1), .IN7(1'b0), .IN8(na3793_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a981_4 ( .OUT(na981_2), .IN1(na1202_1), .IN2(1'b0), .IN3(na1204_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y99     80'h00_0018_00_0040_0A64_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a982_1 ( .OUT(na982_1), .IN1(~na1210_1), .IN2(1'b1), .IN3(na1204_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1214_1), .IN7(~na4328_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x95y100     80'h00_0018_00_0000_0666_5BED
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a984_1 ( .OUT(na984_1), .IN1(na977_1), .IN2(~na4295_2), .IN3(~na4292_2), .IN4(~na3793_2), .IN5(~na977_2), .IN6(na4296_2),
                     .IN7(na987_2), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x96y97     80'h00_0060_00_0000_0C06_FF3D
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a987_4 ( .OUT(na987_2), .IN1(na3790_1), .IN2(~na979_2), .IN3(1'b1), .IN4(na1208_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x94y99     80'h00_0018_00_0000_0666_C606
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a989_1 ( .OUT(na989_1), .IN1(na1210_1), .IN2(na991_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1200_1), .IN6(na3792_2), .IN7(1'b0),
                     .IN8(na992_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y98     80'h00_0018_00_0040_0AE1_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a991_1 ( .OUT(na991_1), .IN1(~na977_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na3793_2), .IN5(1'b1), .IN6(na979_1), .IN7(na4327_2),
                     .IN8(na3793_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y102     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a992_1 ( .OUT(na992_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na979_2), .IN7(1'b1), .IN8(na981_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x100y97     80'h00_0018_00_0000_0C88_95FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a993_1 ( .OUT(na993_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4291_2), .IN6(1'b0), .IN7(~na1212_1), .IN8(~na1208_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y100     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a994_1 ( .OUT(na994_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4288_2), .IN5(~na1202_1), .IN6(1'b0), .IN7(~na1204_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y101     80'h00_0018_00_0040_0AF5_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_1 ( .OUT(na995_1), .IN1(1'b1), .IN2(na984_1), .IN3(na989_1), .IN4(1'b1), .IN5(~na1852_1), .IN6(na3796_1), .IN7(~na4419_2),
                     .IN8(na3800_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y101     80'h00_0018_00_0040_0A7C_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a996_1 ( .OUT(na996_1), .IN1(1'b1), .IN2(na998_1), .IN3(1'b1), .IN4(na997_1), .IN5(na4416_2), .IN6(na979_2), .IN7(~na1013_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x94y102     80'h00_0018_00_0040_0AF5_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a997_1 ( .OUT(na997_1), .IN1(~na1852_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4298_2), .IN5(~na3798_1), .IN6(na4417_2), .IN7(~na989_1),
                     .IN8(na3800_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y102     80'h00_0018_00_0040_0AF5_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a998_1 ( .OUT(na998_1), .IN1(1'b1), .IN2(na984_1), .IN3(1'b1), .IN4(na3800_2), .IN5(~na1852_1), .IN6(na4364_2), .IN7(~na989_1),
                     .IN8(na3800_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x111y102     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_1 ( .OUT(na999_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1000_1), .IN6(1'b0), .IN7(na1004_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y103     80'h00_0018_00_0040_0A74_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1), .IN1(1'b1), .IN2(na998_1), .IN3(1'b1), .IN4(na997_1), .IN5(na3801_1), .IN6(na1001_2), .IN7(~na4300_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x99y102     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1001_4 ( .OUT(na1001_2), .IN1(~na977_1), .IN2(1'b0), .IN3(1'b0), .IN4(na978_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x99y101     80'h00_0060_00_0000_0C06_FFC9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1002_4 ( .OUT(na1002_2), .IN1(na1003_1), .IN2(~na979_1), .IN3(1'b0), .IN4(na978_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x103y101     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_1 ( .OUT(na1003_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1204_1), .IN8(na1206_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y103     80'h00_0018_00_0040_0A7E_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1004_1 ( .OUT(na1004_1), .IN1(1'b1), .IN2(~na976_1), .IN3(na995_1), .IN4(1'b1), .IN5(na4420_2), .IN6(~na1005_2), .IN7(~na4304_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x101y102     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1005_4 ( .OUT(na1005_2), .IN1(na1200_1), .IN2(1'b0), .IN3(~na1006_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x100y101     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1006_1 ( .OUT(na1006_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4293_2), .IN6(~na979_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x101y101     80'h00_0018_00_0000_0C66_6500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1007_1 ( .OUT(na1007_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1202_1), .IN6(1'b0), .IN7(na1204_1), .IN8(na4290_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y101     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1008_1 ( .OUT(na1008_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1010_1), .IN6(na1012_1), .IN7(na1009_1),
                      .IN8(~na1011_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y97     80'h00_0018_00_0040_0AD6_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1), .IN1(1'b1), .IN2(~na976_1), .IN3(1'b1), .IN4(~na997_1), .IN5(na4294_2), .IN6(1'b1), .IN7(~na1013_2),
                      .IN8(na3793_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y99     80'h00_0018_00_0040_0AB5_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_1 ( .OUT(na1010_1), .IN1(1'b1), .IN2(~na998_1), .IN3(na995_1), .IN4(1'b1), .IN5(~na977_1), .IN6(na3804_1), .IN7(1'b1),
                      .IN8(na4290_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y102     80'h00_0018_00_0040_0A76_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1011_1 ( .OUT(na1011_1), .IN1(1'b1), .IN2(na998_1), .IN3(1'b1), .IN4(na997_1), .IN5(na977_1), .IN6(~na4289_2), .IN7(~na4421_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y102     80'h00_0018_00_0040_0A7E_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_1 ( .OUT(na1012_1), .IN1(1'b1), .IN2(~na976_1), .IN3(na995_1), .IN4(1'b1), .IN5(na3806_2), .IN6(~na4301_2), .IN7(~na1013_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x102y101     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1013_4 ( .OUT(na1013_2), .IN1(1'b0), .IN2(na979_2), .IN3(1'b0), .IN4(na3793_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x113y101     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1014_1 ( .OUT(na1014_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1015_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1016_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y103     80'h00_0018_00_0040_0AB7_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1015_1 ( .OUT(na1015_1), .IN1(1'b1), .IN2(na976_1), .IN3(1'b1), .IN4(na997_1), .IN5(~na1200_1), .IN6(~na1005_2), .IN7(1'b1),
                      .IN8(na4303_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y102     80'h00_0018_00_0040_0A7E_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_1 ( .OUT(na1016_1), .IN1(1'b1), .IN2(na998_1), .IN3(na995_1), .IN4(1'b1), .IN5(na4422_2), .IN6(~na1001_2), .IN7(~na4304_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x136y89     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1017_1 ( .OUT(na1017_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3809_2), .IN8(na972_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1017_2 ( .OUT(na1017_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1017_1_i) );
// C_XOR////D      x145y94     80'h40_E818_00_0000_0666_C00A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_1 ( .OUT(na1018_1), .IN1(na1019_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1022_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1018_5 ( .OUT(na1018_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1018_1) );
// C_XOR////      x111y101     80'h00_0018_00_0000_0666_693A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1019_1 ( .OUT(na1019_1), .IN1(na975_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na1016_1), .IN5(~na1015_1), .IN6(na1012_1), .IN7(na996_1),
                      .IN8(na1011_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x100y94     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1022_4 ( .OUT(na1022_2), .IN1(~na1026_1), .IN2(na999_1), .IN3(na1023_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y95     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1023_4 ( .OUT(na1023_2), .IN1(na1010_1), .IN2(~na1025_1), .IN3(na1009_1), .IN4(~na1024_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y98     80'h00_0018_00_0040_0AE8_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1024_1 ( .OUT(na1024_1), .IN1(1'b1), .IN2(~na998_1), .IN3(~na995_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1005_2), .IN7(na4304_2),
                      .IN8(~na3802_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y98     80'h00_0018_00_0040_0AE3_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1), .IN1(1'b1), .IN2(na976_1), .IN3(1'b1), .IN4(~na997_1), .IN5(1'b1), .IN6(~na1001_2), .IN7(na1006_1),
                      .IN8(na3811_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y99     80'h00_0018_00_0000_0C66_5C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1026_1 ( .OUT(na1026_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1028_1), .IN7(~na1027_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y97     80'h00_0018_00_0040_0AB8_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1027_1 ( .OUT(na1027_1), .IN1(1'b1), .IN2(~na998_1), .IN3(1'b1), .IN4(na997_1), .IN5(na1007_1), .IN6(na1001_2), .IN7(1'b0),
                      .IN8(~na3808_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y100     80'h00_0018_00_0040_0AE3_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1), .IN1(1'b1), .IN2(na976_1), .IN3(~na995_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1005_2), .IN7(na4300_2),
                      .IN8(na3813_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x145y88     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1029_1 ( .OUT(na1029_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3814_1), .IN6(na1018_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1029_2 ( .OUT(na1029_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1029_1_i) );
// C_XOR////D      x140y96     80'h40_E818_00_0000_0666_C05C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1), .IN1(1'b0), .IN2(na973_1), .IN3(~na1033_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1031_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1030_5 ( .OUT(na1030_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1030_1) );
// C_XOR////      x114y102     80'h00_0018_00_0000_0C66_5600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1031_1 ( .OUT(na1031_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4308_2), .IN6(na999_1), .IN7(~na1032_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x108y101     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1032_1 ( .OUT(na1032_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na975_2), .IN6(na1028_1), .IN7(~na1027_1),
                      .IN8(na4299_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y101     80'h00_0018_00_0000_0666_9969
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1), .IN1(na975_2), .IN2(~na4305_2), .IN3(na1032_1), .IN4(na1011_1), .IN5(~na1015_1), .IN6(na1012_1),
                      .IN7(na996_1), .IN8(~na1016_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x142y92     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1034_1 ( .OUT(na1034_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4425_2), .IN8(na1030_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1034_2 ( .OUT(na1034_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1034_1_i) );
// C_XOR////D      x142y100     80'h40_E818_00_0000_0666_A03C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_1 ( .OUT(na1035_1), .IN1(1'b0), .IN2(na973_1), .IN3(1'b0), .IN4(~na1036_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1033_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1035_5 ( .OUT(na1035_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1035_1) );
// C_XOR////      x110y100     80'h00_0018_00_0000_0666_AA39
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1036_1 ( .OUT(na1036_1), .IN1(~na1008_1), .IN2(na1028_1), .IN3(1'b0), .IN4(~na1038_1), .IN5(na1039_1), .IN6(1'b0), .IN7(na1027_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y100     80'h00_0018_00_0040_0AD1_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1038_1 ( .OUT(na1038_1), .IN1(1'b1), .IN2(~na976_1), .IN3(~na995_1), .IN4(1'b1), .IN5(~na977_2), .IN6(1'b0), .IN7(na3816_1),
                      .IN8(na4307_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y99     80'h00_0018_00_0040_0ABD_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1), .IN1(1'b1), .IN2(~na998_1), .IN3(1'b1), .IN4(na997_1), .IN5(~na977_1), .IN6(na3817_2), .IN7(1'b1),
                      .IN8(~na4302_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x128y83     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1040_1 ( .OUT(na1040_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3818_1), .IN8(na1035_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1040_2 ( .OUT(na1040_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1040_1_i) );
// C_XOR////D      x135y95     80'h40_E818_00_0000_0666_6003
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1041_1 ( .OUT(na1041_1), .IN1(1'b0), .IN2(~na1042_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1033_1), .IN8(na1036_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1041_5 ( .OUT(na1041_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1041_1) );
// C_///XOR/      x107y98     80'h00_0060_00_0000_0C06_FF96
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1042_4 ( .OUT(na1042_2), .IN1(na1008_1), .IN2(na1025_1), .IN3(~na1032_1), .IN4(na1024_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x137y84     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1044_1 ( .OUT(na1044_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1041_1), .IN6(na3819_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1044_2 ( .OUT(na1044_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1044_1_i) );
// C_XOR////D      x128y91     80'h40_E818_00_0000_0666_A009
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1045_1 ( .OUT(na1045_1), .IN1(~na1026_1), .IN2(na1046_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1047_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1045_5 ( .OUT(na1045_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1045_1) );
// C_XOR////      x107y98     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1046_1 ( .OUT(na1046_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1008_1), .IN6(~na999_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x96y95     80'h00_0018_00_0000_0666_9C96
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1047_1 ( .OUT(na1047_1), .IN1(na1039_1), .IN2(na1028_1), .IN3(~na1027_1), .IN4(na1024_1), .IN5(1'b0), .IN6(na1025_1), .IN7(na1032_1),
                      .IN8(~na1038_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x122y84     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1048_1 ( .OUT(na1048_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1045_1), .IN8(na3820_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1048_2 ( .OUT(na1048_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1048_1_i) );
// C_XOR////D      x134y82     80'h40_E818_00_0000_0666_A0A0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1049_1 ( .OUT(na1049_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1047_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1023_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1049_5 ( .OUT(na1049_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1049_1) );
// C_MX2b/D///      x132y78     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1050_1 ( .OUT(na1050_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4429_2), .IN8(na1049_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1050_2 ( .OUT(na1050_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1050_1_i) );
// C_XOR////D      x138y77     80'h40_E818_00_0000_0666_A030
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_1 ( .OUT(na1051_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(~na1022_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1047_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1051_5 ( .OUT(na1051_2), .CLK(1'b0), .EN(na26_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1051_1) );
// C_MX2b/D///      x131y75     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1052_1 ( .OUT(na1052_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1051_1), .IN8(na3822_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1052_2 ( .OUT(na1052_1), .CLK(1'b0), .EN(na1466_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1052_1_i) );
// C_MX2b/D///      x130y82     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1053_1 ( .OUT(na1053_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na816_1), .IN7(1'b0), .IN8(na3730_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1053_2 ( .OUT(na1053_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1053_1_i) );
// C_MX2b/D///      x123y85     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1054_1 ( .OUT(na1054_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na862_1), .IN7(1'b0), .IN8(na3735_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1054_2 ( .OUT(na1054_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1054_1_i) );
// C_MX2b/D///      x135y83     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_1 ( .OUT(na1055_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na871_1), .IN7(1'b0), .IN8(na4391_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1055_2 ( .OUT(na1055_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1055_1_i) );
// C_MX2b/D///      x135y74     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1056_1 ( .OUT(na1056_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na877_1), .IN7(1'b0), .IN8(na4392_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1056_2 ( .OUT(na1056_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1056_1_i) );
// C_MX2b/D///      x125y78     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1057_1 ( .OUT(na1057_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_1), .IN5(1'b0), .IN6(na4393_2), .IN7(1'b0), .IN8(na883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1057_2 ( .OUT(na1057_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1057_1_i) );
// C_MX2b/D///      x130y76     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1058_1 ( .OUT(na1058_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na887_1), .IN7(1'b0), .IN8(na4394_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1058_2 ( .OUT(na1058_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1058_1_i) );
// C_MX2b/D///      x130y70     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_1 ( .OUT(na1059_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_1), .IN5(1'b0), .IN6(na3742_2), .IN7(1'b0), .IN8(na890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1059_2 ( .OUT(na1059_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1059_1_i) );
// C_MX2b/D///      x131y68     80'h40_E800_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1060_1 ( .OUT(na1060_1_i), .IN1(1'b1), .IN2(~na4175_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na892_1), .IN8(na3743_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1060_2 ( .OUT(na1060_1), .CLK(1'b0), .EN(na1452_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1060_1_i) );
// C_MX2b/D///      x152y96     80'h40_E400_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_1 ( .OUT(na1061_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_1), .IN5(1'b0), .IN6(na3770_1), .IN7(1'b0), .IN8(na895_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1061_2 ( .OUT(na1061_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1061_1_i) );
// C_MX2b/D///      x147y96     80'h40_E400_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1062_1 ( .OUT(na1062_1_i), .IN1(1'b1), .IN2(~na4175_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4285_2), .IN8(na3775_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1062_2 ( .OUT(na1062_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1062_1_i) );
// C_MX2b/D///      x150y96     80'h40_E400_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_1 ( .OUT(na1063_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_1), .IN5(1'b0), .IN6(na3776_2), .IN7(1'b0), .IN8(na949_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1063_2 ( .OUT(na1063_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1063_1_i) );
// C_MX2b/D///      x150y91     80'h40_E400_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_1), .IN5(na955_1), .IN6(1'b0), .IN7(na4410_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1064_2 ( .OUT(na1064_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1064_1_i) );
// C_MX2b/D///      x147y91     80'h40_E400_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1065_1 ( .OUT(na1065_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na25_1), .IN5(na3780_2), .IN6(1'b0), .IN7(na962_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1065_2 ( .OUT(na1065_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1065_1_i) );
// C_MX2b/D///      x150y88     80'h40_E400_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1066_1 ( .OUT(na1066_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na965_1), .IN7(1'b0), .IN8(na3781_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1066_2 ( .OUT(na1066_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1066_1_i) );
// C_MX2b/D///      x137y79     80'h40_E400_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1067_1 ( .OUT(na1067_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na968_1), .IN7(1'b0), .IN8(na3782_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1067_2 ( .OUT(na1067_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1067_1_i) );
// C_MX2b/D///      x144y75     80'h40_E400_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1068_1 ( .OUT(na1068_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_1), .IN5(na970_1), .IN6(1'b0), .IN7(na3783_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1068_2 ( .OUT(na1068_1), .CLK(1'b0), .EN(~na1465_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1068_1_i) );
// C_MX2b/D///      x140y89     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_1 ( .OUT(na1069_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3809_2), .IN8(na972_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1069_2 ( .OUT(na1069_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1069_1_i) );
// C_MX2b/D///      x140y87     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3814_1), .IN6(na1018_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1070_2 ( .OUT(na1070_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1070_1_i) );
// C_MX2b/D///      x143y92     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_1 ( .OUT(na1071_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4425_2), .IN8(na1030_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1071_2 ( .OUT(na1071_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1071_1_i) );
// C_MX2b/D///      x140y85     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1072_1 ( .OUT(na1072_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3818_1), .IN8(na1035_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1072_2 ( .OUT(na1072_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1072_1_i) );
// C_MX2b/D///      x135y87     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1073_1 ( .OUT(na1073_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1041_1), .IN6(na3819_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1073_2 ( .OUT(na1073_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1073_1_i) );
// C_MX2a/D///      x128y85     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1074_1 ( .OUT(na1074_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1045_1), .IN4(na3820_1), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1074_2 ( .OUT(na1074_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1074_1_i) );
// C_MX2b/D///      x140y79     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1075_1 ( .OUT(na1075_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4429_2), .IN8(na1049_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1075_2 ( .OUT(na1075_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1075_1_i) );
// C_MX2b/D///      x128y69     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1076_1 ( .OUT(na1076_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1051_1), .IN8(na3822_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1076_2 ( .OUT(na1076_1), .CLK(1'b0), .EN(na1455_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1076_1_i) );
// C_MX2b/D///      x133y80     80'h40_E400_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1077_1 ( .OUT(na1077_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4389_2), .IN6(na816_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1077_2 ( .OUT(na1077_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1077_1_i) );
// C_MX2b/D///      x125y83     80'h40_E400_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1078_1 ( .OUT(na1078_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4390_2), .IN6(na862_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1078_2 ( .OUT(na1078_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1078_1_i) );
// C_MX2a/D///      x135y81     80'h40_E400_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_1 ( .OUT(na1079_1_i), .IN1(na3736_1), .IN2(na871_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na21_1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1079_2 ( .OUT(na1079_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1079_1_i) );
// C_MX2b/D///      x135y73     80'h40_E400_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1080_1 ( .OUT(na1080_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3739_2), .IN6(na877_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1080_2 ( .OUT(na1080_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1080_1_i) );
// C_MX2a/D///      x124y74     80'h40_E400_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3740_1), .IN4(na883_1), .IN5(~na21_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1081_2 ( .OUT(na1081_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1081_1_i) );
// C_MX2b/D///      x126y73     80'h40_E400_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1082_1 ( .OUT(na1082_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3741_2), .IN6(na887_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1082_2 ( .OUT(na1082_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1082_1_i) );
// C_MX2b/D///      x136y70     80'h40_E400_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_1 ( .OUT(na1083_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4395_2), .IN8(na890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1083_2 ( .OUT(na1083_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1083_1_i) );
// C_MX2b/D///      x133y68     80'h40_E400_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1084_1 ( .OUT(na1084_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na892_1), .IN8(na3743_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1084_2 ( .OUT(na1084_1), .CLK(1'b0), .EN(~na1463_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1084_1_i) );
// C_MX2b/D///      x146y93     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_1 ( .OUT(na1085_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4407_2), .IN8(na895_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1085_2 ( .OUT(na1085_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1085_1_i) );
// C_MX2a/D///      x145y95     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1086_1 ( .OUT(na1086_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na4285_2), .IN4(na3775_1), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1086_2 ( .OUT(na1086_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1086_1_i) );
// C_MX2b/D///      x150y92     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_1 ( .OUT(na1087_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4409_2), .IN8(na949_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1087_2 ( .OUT(na1087_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1087_1_i) );
// C_MX2a/D///      x148y92     80'h40_E800_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1088_1 ( .OUT(na1088_1_i), .IN1(na955_1), .IN2(na3779_1), .IN3(1'b0), .IN4(1'b0), .IN5(na552_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1088_2 ( .OUT(na1088_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1088_1_i) );
// C_MX2b/D///      x146y91     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1089_1 ( .OUT(na1089_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na962_1), .IN8(na4411_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1089_2 ( .OUT(na1089_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1089_1_i) );
// C_MX2b/D///      x148y83     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1090_1 ( .OUT(na1090_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4412_2), .IN6(na965_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1090_2 ( .OUT(na1090_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1090_1_i) );
// C_MX2b/D///      x143y79     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1091_1 ( .OUT(na1091_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4413_2), .IN6(na968_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1091_2 ( .OUT(na1091_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1091_1_i) );
// C_MX2b/D///      x143y75     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1092_1 ( .OUT(na1092_1_i), .IN1(na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na970_1), .IN6(na4414_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1092_2 ( .OUT(na1092_1), .CLK(1'b0), .EN(na1458_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1092_1_i) );
// C_MX2a/D///      x137y89     80'h40_E800_00_0040_0C0A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1093_1 ( .OUT(na1093_1_i), .IN1(1'b0), .IN2(na4423_2), .IN3(1'b0), .IN4(na972_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na25_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1093_2 ( .OUT(na1093_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1093_1_i) );
// C_MX2b/D///      x140y90     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1094_1 ( .OUT(na1094_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_1), .IN5(1'b0), .IN6(na1018_1), .IN7(1'b0), .IN8(na4424_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1094_2 ( .OUT(na1094_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1094_1_i) );
// C_MX2a/D///      x140y91     80'h40_E800_00_0040_0C0A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1095_1 ( .OUT(na1095_1_i), .IN1(1'b0), .IN2(na3815_2), .IN3(1'b0), .IN4(na1030_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na25_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1095_2 ( .OUT(na1095_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1095_1_i) );
// C_MX2b/D///      x137y86     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1096_1 ( .OUT(na1096_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na4426_2), .IN7(1'b0), .IN8(na1035_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1096_2 ( .OUT(na1096_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1096_1_i) );
// C_MX2b/D///      x139y88     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1097_1 ( .OUT(na1097_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na25_1), .IN5(na1041_1), .IN6(1'b0), .IN7(na4427_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1097_2 ( .OUT(na1097_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1097_1_i) );
// C_MX2b/D///      x133y86     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1098_1 ( .OUT(na1098_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_1), .IN5(na4428_2), .IN6(1'b0), .IN7(na1045_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1098_2 ( .OUT(na1098_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1098_1_i) );
// C_MX2b/D///      x136y80     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1099_1 ( .OUT(na1099_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na3821_1), .IN7(1'b0), .IN8(na1049_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1099_2 ( .OUT(na1099_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1099_1_i) );
// C_MX2a/D///      x135y76     80'h40_E800_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1100_1 ( .OUT(na1100_1_i), .IN1(na4430_2), .IN2(1'b0), .IN3(na1051_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na25_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1100_2 ( .OUT(na1100_1), .CLK(1'b0), .EN(na1472_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1100_1_i) );
// C_MX2b/D///      x118y82     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1101_1 ( .OUT(na1101_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na25_2), .IN5(na3871_1), .IN6(1'b0), .IN7(na214_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1101_2 ( .OUT(na1101_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1101_1_i) );
// C_MX2a/D///      x134y78     80'h40_E800_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1102_1 ( .OUT(na1102_1_i), .IN1(na264_1), .IN2(1'b0), .IN3(na3872_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na25_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1102_2 ( .OUT(na1102_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1102_1_i) );
// C_MX2b/D///      x132y81     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1103_1 ( .OUT(na1103_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_2), .IN5(1'b0), .IN6(na3873_2), .IN7(1'b0), .IN8(na277_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1103_2 ( .OUT(na1103_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1103_1_i) );
// C_MX2b/D///      x130y67     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1104_1 ( .OUT(na1104_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na25_2), .IN5(na3874_1), .IN6(1'b0), .IN7(na287_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1104_2 ( .OUT(na1104_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1104_1_i) );
// C_MX2b/D///      x121y71     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1105_1 ( .OUT(na1105_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na25_2), .IN5(na3875_2), .IN6(1'b0), .IN7(na295_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1105_2 ( .OUT(na1105_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1105_1_i) );
// C_MX2b/D///      x126y69     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1106_1 ( .OUT(na1106_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_2), .IN5(na300_1), .IN6(1'b0), .IN7(na3876_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1106_2 ( .OUT(na1106_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1106_1_i) );
// C_MX2a/D///      x129y65     80'h40_E800_00_0040_0C0A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1107_1 ( .OUT(na1107_1_i), .IN1(1'b0), .IN2(na309_1), .IN3(1'b0), .IN4(na3877_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na25_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1107_2 ( .OUT(na1107_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1107_1_i) );
// C_MX2b/D///      x121y65     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1108_1 ( .OUT(na1108_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_2), .IN5(na315_1), .IN6(1'b0), .IN7(na3878_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1108_2 ( .OUT(na1108_1), .CLK(1'b0), .EN(na1469_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1108_1_i) );
// C_MX2a/D///      x130y81     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1109_1 ( .OUT(na1109_1_i), .IN1(na4389_2), .IN2(na816_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1109_2 ( .OUT(na1109_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1109_1_i) );
// C_MX2b/D///      x124y83     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1110_1 ( .OUT(na1110_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4390_2), .IN6(na862_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1110_2 ( .OUT(na1110_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1110_1_i) );
// C_MX2b/D///      x138y83     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_1 ( .OUT(na1111_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3736_1), .IN6(na871_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1111_2 ( .OUT(na1111_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1111_1_i) );
// C_MX2b/D///      x135y75     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1112_1 ( .OUT(na1112_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3739_2), .IN6(na877_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1112_2 ( .OUT(na1112_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1112_1_i) );
// C_MX2b/D///      x123y78     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1113_1 ( .OUT(na1113_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3740_1), .IN8(na883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1113_2 ( .OUT(na1113_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1113_1_i) );
// C_MX2a/D///      x124y75     80'h40_E800_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1114_1 ( .OUT(na1114_1_i), .IN1(na3741_2), .IN2(na887_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na552_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1114_2 ( .OUT(na1114_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1114_1_i) );
// C_MX2b/D///      x130y71     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1115_1 ( .OUT(na1115_1_i), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4395_2), .IN8(na890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1115_2 ( .OUT(na1115_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1115_1_i) );
// C_MX2a/D///      x132y71     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_1 ( .OUT(na1116_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na892_1), .IN4(na3743_2), .IN5(na552_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1116_2 ( .OUT(na1116_1), .CLK(1'b0), .EN(na1462_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1116_1_i) );
// C_MX2b/D///      x146y95     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1117_1 ( .OUT(na1117_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na3770_1), .IN7(1'b0), .IN8(na895_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1117_2 ( .OUT(na1117_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1117_1_i) );
// C_MX2b/D///      x143y98     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1118_1 ( .OUT(na1118_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_1), .IN5(na4408_2), .IN6(1'b0), .IN7(na4285_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1118_2 ( .OUT(na1118_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1118_1_i) );
// C_MX2b/D///      x150y93     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1119_1 ( .OUT(na1119_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na25_1), .IN5(1'b0), .IN6(na3776_2), .IN7(1'b0), .IN8(na949_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1119_2 ( .OUT(na1119_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1119_1_i) );
// C_MX2b/D///      x150y90     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1120_1 ( .OUT(na1120_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na25_1), .IN5(na955_1), .IN6(1'b0), .IN7(na4410_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1120_2 ( .OUT(na1120_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1120_1_i) );
// C_MX2a/D///      x148y89     80'h40_E800_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_1 ( .OUT(na1121_1_i), .IN1(na3780_2), .IN2(1'b0), .IN3(na962_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na25_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1121_2 ( .OUT(na1121_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1121_1_i) );
// C_MX2b/D///      x147y88     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1122_1 ( .OUT(na1122_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_1), .IN5(1'b0), .IN6(na965_1), .IN7(1'b0), .IN8(na3781_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1122_2 ( .OUT(na1122_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1122_1_i) );
// C_MX2a/D///      x137y82     80'h40_E800_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1123_1 ( .OUT(na1123_1_i), .IN1(1'b0), .IN2(na968_1), .IN3(1'b0), .IN4(na3782_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na25_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1123_2 ( .OUT(na1123_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1123_1_i) );
// C_MX2b/D///      x145y78     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1124_1 ( .OUT(na1124_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na25_1), .IN5(na970_1), .IN6(1'b0), .IN7(na3783_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1124_2 ( .OUT(na1124_1), .CLK(1'b0), .EN(na1459_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1124_1_i) );
// C_MX2b/D///      x144y85     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1125_1 ( .OUT(na1125_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3809_2), .IN8(na972_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1125_2 ( .OUT(na1125_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1125_1_i) );
// C_MX2b/D///      x145y87     80'h40_E800_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1126_1 ( .OUT(na1126_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3814_1), .IN6(na1018_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1126_2 ( .OUT(na1126_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1126_1_i) );
// C_MX2b/D///      x143y90     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1127_1 ( .OUT(na1127_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4425_2), .IN8(na1030_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1127_2 ( .OUT(na1127_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1127_1_i) );
// C_MX2a/D///      x141y84     80'h40_E800_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1128_1 ( .OUT(na1128_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3818_1), .IN4(na1035_1), .IN5(na21_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1128_2 ( .OUT(na1128_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1128_1_i) );
// C_MX2b/D///      x135y88     80'h40_E800_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1041_1), .IN6(na3819_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1129_2 ( .OUT(na1129_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1129_1_i) );
// C_MX2a/D///      x128y84     80'h40_E800_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1130_1 ( .OUT(na1130_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1045_1), .IN4(na3820_1), .IN5(~na21_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1130_2 ( .OUT(na1130_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1130_1_i) );
// C_MX2b/D///      x140y75     80'h40_E800_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4429_2), .IN8(na1049_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1131_2 ( .OUT(na1131_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1131_1_i) );
// C_MX2b/D///      x136y76     80'h40_E800_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1132_1 ( .OUT(na1132_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1051_1), .IN8(na3822_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1132_2 ( .OUT(na1132_1), .CLK(1'b0), .EN(na1460_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1132_1_i) );
// C_MX2b/D///      x126y80     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1133_1 ( .OUT(na1133_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1451_2), .IN5(na3871_1), .IN6(1'b0), .IN7(na214_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1133_2 ( .OUT(na1133_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1133_1_i) );
// C_MX2b/D///      x137y74     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(na264_1), .IN6(1'b0), .IN7(na3872_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1134_2 ( .OUT(na1134_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1134_1_i) );
// C_MX2a/D///      x139y78     80'h40_E800_00_0040_0C0A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1_i), .IN1(1'b0), .IN2(na3873_2), .IN3(1'b0), .IN4(na277_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1135_2 ( .OUT(na1135_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1135_1_i) );
// C_MX2b/D///      x136y65     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1136_1 ( .OUT(na1136_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1451_2), .IN5(na3874_1), .IN6(1'b0), .IN7(na287_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1136_2 ( .OUT(na1136_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1136_1_i) );
// C_MX2a/D///      x131y66     80'h40_E800_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1_i), .IN1(na3875_2), .IN2(1'b0), .IN3(na295_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1137_2 ( .OUT(na1137_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1137_1_i) );
// C_MX2b/D///      x123y70     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1138_1 ( .OUT(na1138_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(na300_1), .IN6(1'b0), .IN7(na3876_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1138_2 ( .OUT(na1138_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1138_1_i) );
// C_MX2b/D///      x126y63     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(na309_1), .IN7(1'b0), .IN8(na3877_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1139_2 ( .OUT(na1139_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1139_1_i) );
// C_MX2b/D///      x124y62     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1451_2), .IN5(na315_1), .IN6(1'b0), .IN7(na3878_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1140_2 ( .OUT(na1140_1), .CLK(1'b0), .EN(na1471_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1140_1_i) );
// C_MX2b////D      x132y77     80'h40_E818_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1142_1), .IN4(1'b1), .IN5(na3871_1), .IN6(1'b0), .IN7(na214_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1141_5 ( .OUT(na1141_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1141_1) );
// C_AND////      x138y71     80'h00_0018_00_0000_0C88_82FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1142_1 ( .OUT(na1142_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1335_1), .IN6(~na1333_2), .IN7(na4342_2),
                      .IN8(na1336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////D      x139y74     80'h40_E818_00_0040_0C05_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1143_1 ( .OUT(na1143_1), .IN1(na264_1), .IN2(1'b0), .IN3(na3872_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1142_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1143_5 ( .OUT(na1143_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1143_1) );
// C_MX2a////D      x140y80     80'h40_E818_00_0040_0C0A_5F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1144_1 ( .OUT(na1144_1), .IN1(1'b0), .IN2(na3873_2), .IN3(1'b0), .IN4(na277_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1142_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1144_5 ( .OUT(na1144_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1144_1) );
// C_MX2b////D      x138y66     80'h40_E818_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_1 ( .OUT(na1145_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1142_1), .IN4(1'b1), .IN5(na3874_1), .IN6(1'b0), .IN7(na287_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1145_5 ( .OUT(na1145_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1145_1) );
// C_MX2b////D      x140y67     80'h40_E818_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1146_1 ( .OUT(na1146_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1142_1), .IN4(1'b1), .IN5(na3875_2), .IN6(1'b0), .IN7(na295_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1146_5 ( .OUT(na1146_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1146_1) );
// C_MX2a////D      x133y66     80'h40_E818_00_0040_0C05_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1), .IN1(na300_1), .IN2(1'b0), .IN3(na3876_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1142_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1147_5 ( .OUT(na1147_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1147_1) );
// C_MX2b////D      x127y64     80'h40_E818_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1148_1 ( .OUT(na1148_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1142_1), .IN4(1'b1), .IN5(1'b0), .IN6(na309_1), .IN7(1'b0), .IN8(na3877_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1148_5 ( .OUT(na1148_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1148_1) );
// C_MX2a////D      x124y63     80'h40_E818_00_0040_0C05_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1149_1 ( .OUT(na1149_1), .IN1(na315_1), .IN2(1'b0), .IN3(na3878_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1142_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1149_5 ( .OUT(na1149_2), .CLK(1'b0), .EN(na349_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1149_1) );
// C_///AND/D      x149y61     80'h40_F800_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1150_4 ( .OUT(na1150_2_i), .IN1(na1319_1), .IN2(1'b1), .IN3(1'b1), .IN4(na547_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1150_5 ( .OUT(na1150_2), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1150_2_i) );
// C_MX2b/D///      x89y96     80'h40_EC00_00_0040_0A32_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_1 ( .OUT(na1151_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3871_1), .IN6(~na1153_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1151_2 ( .OUT(na1151_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1151_1_i) );
// C_MX2b////      x97y88     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1153_1 ( .OUT(na1153_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na584_1), .IN6(~na551_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x89y91     80'h40_EC00_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_1 ( .OUT(na1154_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3872_1), .IN8(~na1155_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1154_2 ( .OUT(na1154_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1154_1_i) );
// C_MX2b////      x112y88     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_1 ( .OUT(na1155_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na553_1), .IN6(~na585_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x90y94     80'h40_EC00_00_0040_0C13_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1156_1 ( .OUT(na1156_1_i), .IN1(~na1157_1), .IN2(na3873_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3871_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1156_2 ( .OUT(na1156_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1156_1_i) );
// C_MX2b////      x105y89     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_1 ( .OUT(na1157_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na586_1), .IN6(~na554_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x98y87     80'h40_EC00_00_0040_0C23_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1158_1 ( .OUT(na1158_1_i), .IN1(na3874_1), .IN2(~na1159_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3871_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1158_2 ( .OUT(na1158_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1158_1_i) );
// C_MX2b////      x107y82     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1159_1 ( .OUT(na1159_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na555_1), .IN6(~na587_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x88y93     80'h40_EC00_00_0040_0A32_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1160_1 ( .OUT(na1160_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3875_2), .IN6(~na1161_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1160_2 ( .OUT(na1160_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1160_1_i) );
// C_MX2b////      x99y88     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_1 ( .OUT(na1161_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4203_2), .IN8(~na588_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x87y91     80'h40_EC00_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1162_1 ( .OUT(na1162_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3876_2), .IN8(~na1163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1162_2 ( .OUT(na1162_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1162_1_i) );
// C_MX2a////      x94y86     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_1 ( .OUT(na1163_1), .IN1(~na589_1), .IN2(~na557_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1333_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x88y88     80'h40_EC00_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1164_1 ( .OUT(na1164_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1165_1),
                      .IN8(na3877_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1164_2 ( .OUT(na1164_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1164_1_i) );
// C_MX2a////      x94y79     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1), .IN1(~na558_1), .IN2(~na590_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1333_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x87y88     80'h40_EC00_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1166_1 ( .OUT(na1166_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3878_2), .IN8(~na1167_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1166_2 ( .OUT(na1166_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1166_1_i) );
// C_MX2b////      x98y76     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1167_1 ( .OUT(na1167_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na559_1), .IN8(~na591_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x89y99     80'h40_EC00_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1169_1),
                      .IN8(na3730_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1168_2 ( .OUT(na1168_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1168_1_i) );
// C_MX2b////      x96y91     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1169_1 ( .OUT(na1169_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na560_1), .IN6(~na4221_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x91y97     80'h40_EC00_00_0040_0C4C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_1 ( .OUT(na1170_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1171_1), .IN4(na3735_1), .IN5(~na3871_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1170_2 ( .OUT(na1170_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1170_1_i) );
// C_MX2b////      x106y89     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_1 ( .OUT(na1171_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na561_1), .IN6(~na593_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x92y100     80'h40_EC00_00_0040_0C23_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1172_1 ( .OUT(na1172_1_i), .IN1(na3736_1), .IN2(~na1173_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3871_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1172_2 ( .OUT(na1172_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1172_1_i) );
// C_MX2b////      x103y88     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_1 ( .OUT(na1173_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na594_1), .IN6(~na562_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x91y94     80'h40_EC00_00_0040_0A32_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1174_1 ( .OUT(na1174_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3739_2), .IN6(~na1175_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1174_2 ( .OUT(na1174_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1174_1_i) );
// C_MX2b////      x109y78     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1175_1 ( .OUT(na1175_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na563_1), .IN6(~na595_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x90y95     80'h40_EC00_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1176_1 ( .OUT(na1176_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3740_1), .IN8(~na1177_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1176_2 ( .OUT(na1176_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1176_1_i) );
// C_MX2a////      x102y84     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1177_1 ( .OUT(na1177_1), .IN1(~na564_1), .IN2(~na596_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1333_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x93y99     80'h40_EC00_00_0040_0A32_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1178_1 ( .OUT(na1178_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3741_2), .IN6(~na1179_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1178_2 ( .OUT(na1178_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1178_1_i) );
// C_MX2a////      x93y86     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1179_1 ( .OUT(na1179_1), .IN1(~na597_1), .IN2(~na4204_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1333_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x89y90     80'h40_EC00_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1180_1 ( .OUT(na1180_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1181_1), .IN6(na3742_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1180_2 ( .OUT(na1180_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1180_1_i) );
// C_MX2b////      x93y77     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1181_1 ( .OUT(na1181_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na598_1), .IN8(~na4206_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x92y93     80'h40_EC00_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1182_1 ( .OUT(na1182_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1183_1),
                      .IN8(na3743_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1182_2 ( .OUT(na1182_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1182_1_i) );
// C_MX2b////      x96y75     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1183_1 ( .OUT(na1183_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4223_2), .IN8(~na567_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x120y95     80'h40_EC00_00_0040_0C13_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1184_1 ( .OUT(na1184_1_i), .IN1(~na1185_1), .IN2(na3770_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3871_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1184_2 ( .OUT(na1184_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1184_1_i) );
// C_MX2b////      x129y95     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1185_1 ( .OUT(na1185_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na568_1), .IN6(~na600_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x124y100     80'h40_EC00_00_0040_0C4C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1186_1 ( .OUT(na1186_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1187_1), .IN4(na3775_1), .IN5(~na3871_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1186_2 ( .OUT(na1186_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1186_1_i) );
// C_MX2b////      x132y99     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1187_1 ( .OUT(na1187_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na569_1), .IN6(~na601_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x119y100     80'h40_EC00_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1188_1 ( .OUT(na1188_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1189_1), .IN6(na3776_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1188_2 ( .OUT(na1188_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1188_1_i) );
// C_MX2b////      x129y97     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1189_1 ( .OUT(na1189_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na602_1), .IN6(~na4208_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x129y93     80'h40_EC00_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1190_1 ( .OUT(na1190_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1191_1), .IN6(na3779_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1190_2 ( .OUT(na1190_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1190_1_i) );
// C_MX2a////      x127y87     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1191_1 ( .OUT(na1191_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na603_1), .IN4(~na4210_2), .IN5(1'b1), .IN6(~na1333_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x115y101     80'h40_EC00_00_0040_0A32_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1192_1 ( .OUT(na1192_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3780_2), .IN6(~na1193_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1192_2 ( .OUT(na1192_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1192_1_i) );
// C_MX2a////      x121y88     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1193_1 ( .OUT(na1193_1), .IN1(~na572_1), .IN2(~na604_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1333_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x112y94     80'h40_EC00_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1194_1 ( .OUT(na1194_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1195_1),
                      .IN8(na3781_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1194_2 ( .OUT(na1194_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1194_1_i) );
// C_MX2b////      x118y85     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1195_1 ( .OUT(na1195_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na605_1), .IN6(~na573_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x127y86     80'h40_EC00_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1196_1 ( .OUT(na1196_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1197_1),
                      .IN8(na3782_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1196_2 ( .OUT(na1196_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1196_1_i) );
// C_MX2b////      x112y75     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1197_1 ( .OUT(na1197_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na606_1), .IN6(~na4211_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x114y87     80'h40_EC00_00_0040_0C8C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1198_1 ( .OUT(na1198_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3783_1), .IN4(~na1199_1), .IN5(na3871_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1198_2 ( .OUT(na1198_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1198_1_i) );
// C_MX2b////      x120y78     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_1 ( .OUT(na1199_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na575_1), .IN6(~na607_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x111y99     80'h40_EC00_00_0040_0C8C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1200_1 ( .OUT(na1200_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3809_2), .IN4(~na1201_1), .IN5(na3871_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1200_2 ( .OUT(na1200_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1200_1_i) );
// C_MX2b////      x110y92     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1201_1 ( .OUT(na1201_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na576_1), .IN6(~na608_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x109y97     80'h40_EC00_00_0040_0A32_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1202_1 ( .OUT(na1202_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3814_1), .IN6(~na1203_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1202_2 ( .OUT(na1202_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1202_1_i) );
// C_MX2b////      x117y86     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1203_1 ( .OUT(na1203_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na4214_2), .IN6(~na609_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x110y101     80'h40_EC00_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1204_1 ( .OUT(na1204_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1205_1), .IN6(na3815_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1204_2 ( .OUT(na1204_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1204_1_i) );
// C_MX2a////      x115y93     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1205_1 ( .OUT(na1205_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na578_1), .IN4(~na610_1), .IN5(1'b1), .IN6(na1333_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x116y100     80'h40_EC00_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1206_1 ( .OUT(na1206_1_i), .IN1(na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3818_1), .IN8(~na1207_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1206_2 ( .OUT(na1206_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1206_1_i) );
// C_MX2a////      x112y90     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1207_1 ( .OUT(na1207_1), .IN1(~na579_1), .IN2(~na611_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1333_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x112y100     80'h40_EC00_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1208_1 ( .OUT(na1208_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1209_1), .IN6(na3819_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1208_2 ( .OUT(na1208_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1208_1_i) );
// C_MX2b////      x109y89     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1209_1 ( .OUT(na1209_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na580_1), .IN6(~na612_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x105y101     80'h40_EC00_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1210_1 ( .OUT(na1210_1_i), .IN1(~na3871_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1211_1),
                      .IN8(na3820_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1210_2 ( .OUT(na1210_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1210_1_i) );
// C_MX2b////      x102y85     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1211_1 ( .OUT(na1211_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na613_1), .IN6(~na4217_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x98y95     80'h40_EC00_00_0040_0C13_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1212_1 ( .OUT(na1212_1_i), .IN1(~na1213_1), .IN2(na3821_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3871_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1212_2 ( .OUT(na1212_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1212_1_i) );
// C_MX2b////      x107y79     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1213_1 ( .OUT(na1213_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na614_1), .IN6(~na4219_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x109y98     80'h40_EC00_00_0040_0C4C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1214_1 ( .OUT(na1214_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1215_1), .IN4(na3822_2), .IN5(~na3871_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1214_2 ( .OUT(na1214_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1214_1_i) );
// C_MX2b////      x106y79     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1215_1 ( .OUT(na1215_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na583_1), .IN8(~na615_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x147y64     80'h40_F800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1216_4 ( .OUT(na1216_2_i), .IN1(1'b1), .IN2(na1912_1), .IN3(1'b1), .IN4(~na547_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1216_5 ( .OUT(na1216_2), .CLK(1'b0), .EN(na1396_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1216_2_i) );
// C_AND/D//AND/D      x152y63     80'h40_F800_80_0000_0C88_3C1F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1217_1 ( .OUT(na1217_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1912_2), .IN7(1'b1), .IN8(~na547_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1217_2 ( .OUT(na1217_1), .CLK(1'b0), .EN(na1396_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1217_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1217_4 ( .OUT(na1217_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1217_2), .IN4(~na547_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1217_5 ( .OUT(na1217_2), .CLK(1'b0), .EN(na1396_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1217_2_i) );
// C_OR/D///      x150y78     80'h40_E800_00_0000_0EEE_B03D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1219_1 ( .OUT(na1219_1_i), .IN1(~na3952_1), .IN2(na3970_1), .IN3(1'b0), .IN4(~na3967_2), .IN5(1'b0), .IN6(1'b0), .IN7(na3968_1),
                      .IN8(~na3967_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1219_2 ( .OUT(na1219_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1219_1_i) );
// C_///AND/      x154y86     80'h00_0060_00_0000_0C08_FFC8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1222_4 ( .OUT(na1222_2), .IN1(na10_1), .IN2(na12_2), .IN3(1'b1), .IN4(na1223_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y76     80'h00_0018_00_0000_0C88_C1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1223_1 ( .OUT(na1223_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10_2), .IN6(~na12_1), .IN7(1'b1), .IN8(na9_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x154y74     80'h00_0078_00_0000_0C88_AAC8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1224_1 ( .OUT(na1224_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na546_2), .IN6(1'b1), .IN7(na1225_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1224_4 ( .OUT(na1224_2), .IN1(na10_1), .IN2(na12_2), .IN3(1'b1), .IN4(na1239_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x154y75     80'h00_0060_00_0000_0C08_FFC2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1225_4 ( .OUT(na1225_2), .IN1(na10_2), .IN2(~na12_1), .IN3(1'b1), .IN4(na9_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y67     80'h00_0018_00_0000_0C88_31FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1228_1 ( .OUT(na1228_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10_2), .IN6(~na12_1), .IN7(1'b1), .IN8(~na9_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x153y72     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1229_1 ( .OUT(na1229_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(na12_2), .IN7(na1228_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x154y86     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1230_1 ( .OUT(na1230_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3958_1), .IN6(na3297_1), .IN7(1'b0), .IN8(na4167_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y83     80'h00_0018_00_0000_0888_8811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1233_1 ( .OUT(na1233_1), .IN1(~na3962_2), .IN2(~na3960_2), .IN3(~na3966_1), .IN4(~na3964_2), .IN5(na3963_1), .IN6(na3961_1),
                      .IN7(na3965_1), .IN8(na3959_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x152y76     80'h00_0078_00_0000_0C88_A2CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1235_1 ( .OUT(na1235_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(~na12_2), .IN7(na1225_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1235_4 ( .OUT(na1235_2), .IN1(na546_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1239_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x153y77     80'h00_0078_00_0000_0C88_A4A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1236_1 ( .OUT(na1236_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10_1), .IN6(na12_2), .IN7(na1225_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1236_4 ( .OUT(na1236_2), .IN1(na10_1), .IN2(na12_2), .IN3(na1225_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x154y67     80'h00_0060_00_0000_0C08_FFC2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1238_4 ( .OUT(na1238_2), .IN1(na10_1), .IN2(~na12_2), .IN3(1'b1), .IN4(na1239_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y72     80'h00_0018_00_0000_0C88_32FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_1 ( .OUT(na1239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_2), .IN6(~na12_1), .IN7(1'b1), .IN8(~na9_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x153y73     80'h00_0078_00_0000_0C88_A4CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1243_1 ( .OUT(na1243_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10_1), .IN6(na12_2), .IN7(na1228_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1243_4 ( .OUT(na1243_2), .IN1(na546_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1223_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x151y67     80'h00_0078_00_0000_0C88_AAA2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1245_1 ( .OUT(na1245_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na546_2), .IN6(1'b1), .IN7(na1228_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1245_4 ( .OUT(na1245_2), .IN1(na10_1), .IN2(~na12_2), .IN3(na1228_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x152y65     80'h00_0060_00_0000_0C08_FFC4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1246_4 ( .OUT(na1246_2), .IN1(~na10_1), .IN2(na12_2), .IN3(1'b1), .IN4(na1239_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x153y80     80'h00_0078_00_0000_0C88_C2C4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1251_1 ( .OUT(na1251_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(~na12_2), .IN7(1'b1), .IN8(na1223_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1251_4 ( .OUT(na1251_2), .IN1(~na10_1), .IN2(na12_2), .IN3(1'b1), .IN4(na1223_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x153y85     80'h40_E800_00_0000_0EEE_E07C
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1253_1 ( .OUT(na1253_1_i), .IN1(1'b0), .IN2(na3985_1), .IN3(~na3984_2), .IN4(~na3971_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3983_1),
                      .IN8(na1263_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1253_2 ( .OUT(na1253_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1253_1_i) );
// C_///ORAND/      x150y81     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1258_4 ( .OUT(na1258_2), .IN1(~na1078_1), .IN2(~na4337_2), .IN3(~na1110_1), .IN4(~na1224_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x146y78     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1259_1 ( .OUT(na1259_1), .IN1(~na1245_1), .IN2(~na1134_1), .IN3(~na1070_1), .IN4(~na1235_1), .IN5(~na1245_2), .IN6(~na1143_2),
                      .IN7(~na870_1), .IN8(~na1235_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y92     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1263_1 ( .OUT(na1263_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1062_1), .IN7(1'b1), .IN8(na4338_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*/D///      x153y82     80'h40_E800_00_0000_0788_8821
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1265_1 ( .OUT(na1265_1_i), .IN1(~na3987_2), .IN2(~na3989_2), .IN3(na1271_1), .IN4(~na3991_2), .IN5(na1270_1), .IN6(na3986_1),
                      .IN7(na3988_1), .IN8(na3990_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1265_2 ( .OUT(na1265_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1265_1_i) );
// C_ORAND////      x151y87     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1270_1 ( .OUT(na1270_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1236_2), .IN6(~na1127_1), .IN7(~na4310_2),
                      .IN8(~na1224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y79     80'h00_0018_00_0000_0888_8811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_1 ( .OUT(na1271_1), .IN1(~na3999_2), .IN2(~na4001_2), .IN3(~na3997_1), .IN4(~na3995_1), .IN5(na3994_1), .IN6(na3996_2),
                      .IN7(na3998_2), .IN8(na4000_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x151y70     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1277_1 ( .OUT(na1277_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1229_1), .IN7(na1104_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1277_4 ( .OUT(na1277_2), .IN1(na1243_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x152y75     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1280_1 ( .OUT(na1280_1), .IN1(~na1236_1), .IN2(~na1096_1), .IN3(~na1136_1), .IN4(~na4336_2), .IN5(~na1236_2), .IN6(~na1128_1),
                      .IN7(~na4264_2), .IN8(~na1235_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x147y77     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1283_1 ( .OUT(na1283_1), .IN1(~na1080_1), .IN2(~na4337_2), .IN3(~na1040_1), .IN4(~na1224_1), .IN5(~na1112_1), .IN6(~na4330_2),
                      .IN7(~na1072_1), .IN8(~na1235_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x149y70     80'h40_E800_00_0000_0EEE_5CD5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1286_1 ( .OUT(na1286_1_i), .IN1(~na4013_1), .IN2(1'b0), .IN3(~na4025_2), .IN4(na4028_2), .IN5(1'b0), .IN6(na4026_1), .IN7(~na4025_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1286_2 ( .OUT(na1286_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1286_1_i) );
// C_AND////      x147y76     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_1 ( .OUT(na1289_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1113_1), .IN7(1'b1), .IN8(na1224_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x153y89     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1291_1 ( .OUT(na1291_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1236_2), .IN6(~na1129_1), .IN7(~na1121_1),
                      .IN8(~na1222_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1291_4 ( .OUT(na1291_2), .IN1(~na1065_1), .IN2(~na1251_1), .IN3(~na1089_1), .IN4(~na4340_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x146y79     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1293_4 ( .OUT(na1293_2), .IN1(~na1073_1), .IN2(~na4331_2), .IN3(~na886_1), .IN4(~na1235_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x145y74     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1294_1 ( .OUT(na1294_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1105_1), .IN6(~na1229_1), .IN7(~na1246_2),
                      .IN8(~na1081_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x144y71     80'h40_E800_00_0000_0EEE_A5D5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1297_1 ( .OUT(na1297_1_i), .IN1(~na4041_2), .IN2(1'b0), .IN3(~na4029_1), .IN4(na4044_2), .IN5(~na4041_1), .IN6(1'b0), .IN7(na4042_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1297_2 ( .OUT(na1297_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1297_1_i) );
// C_///ORAND/      x151y84     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1302_4 ( .OUT(na1302_2), .IN1(~na1236_1), .IN2(~na1098_1), .IN3(~na1074_1), .IN4(~na1235_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x149y75     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1303_1 ( .OUT(na1303_1), .IN1(~na1243_1), .IN2(~na2923_1), .IN3(~na4265_2), .IN4(~na1235_2), .IN5(~na1243_2), .IN6(~na967_1),
                      .IN7(~na4312_2), .IN8(~na1224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x138y67     80'h40_E800_00_0000_0EEE_3A3D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_1 ( .OUT(na1308_1_i), .IN1(~na4045_1), .IN2(na4060_1), .IN3(1'b0), .IN4(~na4057_2), .IN5(na4058_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(~na4057_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1308_2 ( .OUT(na1308_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1308_1_i) );
// C_AND////      x151y65     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1310_1 ( .OUT(na1310_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2924_2), .IN6(1'b1), .IN7(1'b1), .IN8(na4335_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x152y74     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1067_1), .IN6(~na1251_1), .IN7(~na4313_2),
                      .IN8(~na1224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1313_4 ( .OUT(na1313_2), .IN1(~na1243_2), .IN2(~na969_1), .IN3(~na1238_2), .IN4(~na1059_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x150y75     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1315_1 ( .OUT(na1315_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1091_1), .IN6(~na1251_2), .IN7(~na4266_2),
                      .IN8(~na1235_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x145y74     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1316_4 ( .OUT(na1316_2), .IN1(~na1107_1), .IN2(~na1229_1), .IN3(~na1246_2), .IN4(~na1083_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x145y67     80'h40_E800_00_0000_0EEE_C5C7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1319_1 ( .OUT(na1319_1_i), .IN1(~na4072_2), .IN2(~na4061_1), .IN3(1'b0), .IN4(na4075_1), .IN5(~na4072_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na4073_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1319_2 ( .OUT(na1319_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1319_1_i) );
// C_AND///AND/      x152y69     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_1 ( .OUT(na1323_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1052_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1224_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1323_4 ( .OUT(na1323_2), .IN1(na1243_2), .IN2(na971_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x148y70     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_1 ( .OUT(na1325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4334_2), .IN6(~na1060_1), .IN7(~na4267_2),
                      .IN8(~na1235_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x149y72     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1326_1 ( .OUT(na1326_1), .IN1(~na1092_1), .IN2(~na1251_2), .IN3(~na1068_1), .IN4(~na4339_2), .IN5(~na1243_1), .IN6(~na2925_1),
                      .IN7(~na1116_1), .IN8(~na1224_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x121y67     80'h40_EC00_00_0040_0C9C_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1331_1 ( .OUT(na1331_1_i), .IN1(1'b1), .IN2(1'b0), .IN3(na4076_2), .IN4(~na1332_1), .IN5(na1331_1), .IN6(1'b1), .IN7(na4365_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1331_2 ( .OUT(na1331_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1331_1_i) );
// C_MX4a/DST///      x122y68     80'h60_BC00_00_0040_0C6E_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1332_1 ( .OUT(na1332_1_i), .IN1(1'b0), .IN2(~na1859_1), .IN3(~na4077_1), .IN4(na4366_2), .IN5(na1331_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1332_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0000)) 
           _a1332_2 ( .OUT(na1332_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1332_1_i) );
// C_AND////D      x119y78     80'h40_E418_00_0000_0888_F35F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1142_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1333_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1333_5 ( .OUT(na1333_2), .CLK(1'b0), .EN(~na25_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1333_1) );
// C_AND/D//AND/D      x135y67     80'h40_E400_80_0000_0C88_2F2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1335_1 ( .OUT(na1335_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1883_2), .IN8(~na4314_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1335_2 ( .OUT(na1335_1), .CLK(1'b0), .EN(~na25_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1335_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1335_4 ( .OUT(na1335_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1883_1), .IN4(~na4314_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1335_5 ( .OUT(na1335_2), .CLK(1'b0), .EN(~na25_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1335_2_i) );
// C_///AND/D      x138y64     80'h40_E400_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1336_4 ( .OUT(na1336_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1142_1), .IN4(na1885_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1336_5 ( .OUT(na1336_2), .CLK(1'b0), .EN(~na25_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1336_2_i) );
// C_AND/D///      x87y74     80'h40_EC00_00_0000_0888_8CA2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1337_1 ( .OUT(na1337_1_i), .IN1(na1339_1), .IN2(~na4367_2), .IN3(na1343_1), .IN4(1'b1), .IN5(1'b1), .IN6(na1361_1), .IN7(na1343_2),
                      .IN8(na1345_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1337_2 ( .OUT(na1337_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1337_1_i) );
// C_///AND/      x80y70     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1338_4 ( .OUT(na1338_2), .IN1(na1339_1), .IN2(na4343_2), .IN3(na1343_2), .IN4(na1345_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y59     80'h00_0018_00_0000_0888_8441
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1339_1 ( .OUT(na1339_1), .IN1(~na1358_1), .IN2(~na1355_1), .IN3(~na1359_1), .IN4(na1342_1), .IN5(~na1358_2), .IN6(na1355_2),
                      .IN7(na1359_2), .IN8(na1356_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y64     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1342_1 ( .OUT(na1342_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1351_1), .IN6(~na1353_2), .IN7(~na1357_2),
                      .IN8(~na1346_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x82y65     80'h40_E800_80_0000_0C88_1F3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1343_1 ( .OUT(na1343_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1343_1), .IN8(~na4078_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1343_2 ( .OUT(na1343_1), .CLK(1'b0), .EN(na1448_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1343_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1343_4 ( .OUT(na1343_2_i), .IN1(na1898_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4078_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1343_5 ( .OUT(na1343_2), .CLK(1'b0), .EN(na1448_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1343_2_i) );
// C_AND/D///      x82y68     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1898_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na4078_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1345_2 ( .OUT(na1345_1), .CLK(1'b0), .EN(na1448_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1345_1_i) );
// C_AND/D///      x80y60     80'h40_E400_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1346_1 ( .OUT(na1346_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1347_1), .IN8(~na1346_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1346_2 ( .OUT(na1346_1), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1346_1_i) );
// C_MX2b////      x80y65     80'h00_0018_00_0040_0A32_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1347_1 ( .OUT(na1347_1), .IN1(1'b1), .IN2(~na1361_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1339_1), .IN6(~na4081_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y62     80'h00_0018_00_0000_0888_1441
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1348_1 ( .OUT(na1348_1), .IN1(~na1358_1), .IN2(~na1355_2), .IN3(~na1359_1), .IN4(na1350_2), .IN5(~na1358_2), .IN6(na1355_1),
                      .IN7(~na1359_2), .IN8(~na1356_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x80y64     80'h00_0060_00_0000_0C08_FF48
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1350_4 ( .OUT(na1350_2), .IN1(na1351_1), .IN2(na1353_2), .IN3(~na1357_2), .IN4(na1346_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x81y61     80'h40_E400_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_1 ( .OUT(na1351_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1888_1), .IN6(1'b1), .IN7(~na1347_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1351_2 ( .OUT(na1351_1), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1351_1_i) );
// C_///AND/D      x81y62     80'h40_E400_80_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1353_4 ( .OUT(na1353_2_i), .IN1(1'b1), .IN2(na1890_1), .IN3(~na1347_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1353_5 ( .OUT(na1353_2), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1353_2_i) );
// C_AND/D//AND/D      x81y64     80'h40_E400_80_0000_0C88_5A5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1355_1 ( .OUT(na1355_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1892_1), .IN6(1'b1), .IN7(~na1347_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1355_2 ( .OUT(na1355_1), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1355_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1355_4 ( .OUT(na1355_2_i), .IN1(na1888_2), .IN2(1'b1), .IN3(~na1347_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1355_5 ( .OUT(na1355_2), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1355_2_i) );
// C_///AND/D      x88y64     80'h40_E400_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1356_4 ( .OUT(na1356_2_i), .IN1(na1892_2), .IN2(1'b1), .IN3(~na1347_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1356_5 ( .OUT(na1356_2), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1356_2_i) );
// C_///AND/D      x82y61     80'h40_E400_80_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1357_4 ( .OUT(na1357_2_i), .IN1(1'b1), .IN2(na1894_1), .IN3(~na1347_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1357_5 ( .OUT(na1357_2), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1357_2_i) );
// C_AND/D//AND/D      x83y61     80'h40_E400_80_0000_0C88_5C5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1358_1 ( .OUT(na1358_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1894_2), .IN7(~na1347_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1358_2 ( .OUT(na1358_1), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1358_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1358_4 ( .OUT(na1358_2_i), .IN1(na1896_2), .IN2(1'b1), .IN3(~na1347_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1358_5 ( .OUT(na1358_2), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1358_2_i) );
// C_AND/D//AND/D      x82y63     80'h40_E400_80_0000_0C88_5A5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_1 ( .OUT(na1359_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1896_1), .IN6(1'b1), .IN7(~na1347_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1359_2 ( .OUT(na1359_1), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1359_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1359_4 ( .OUT(na1359_2_i), .IN1(1'b1), .IN2(na1890_2), .IN3(~na1347_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1359_5 ( .OUT(na1359_2), .CLK(1'b0), .EN(~na1449_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1359_2_i) );
// C_XOR/D///      x81y60     80'h40_E800_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1361_1 ( .OUT(na1361_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1361_1), .IN7(na3196_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1361_2 ( .OUT(na1361_1), .CLK(1'b0), .EN(na1397_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1361_1_i) );
// C_MX4a/DST///      x154y58     80'h60_BC00_00_0040_0C92_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1362_1 ( .OUT(na1362_1_i), .IN1(1'b1), .IN2(na1363_1), .IN3(1'b0), .IN4(1'b1), .IN5(~na3235_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1386_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0000)) 
           _a1362_2 ( .OUT(na1362_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1362_1_i) );
// C_MX2b/D///      x153y62     80'h40_F800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_1 ( .OUT(na1363_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na547_1), .IN5(1'b0), .IN6(na1364_1), .IN7(1'b0), .IN8(na1219_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1363_2 ( .OUT(na1363_1), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1363_1_i) );
// C_MX2b/D///      x153y64     80'h40_F800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na547_1), .IN5(na1253_1), .IN6(1'b0), .IN7(na1365_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1364_2 ( .OUT(na1364_1), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1364_1_i) );
// C_MX2b/D///      x154y63     80'h40_F800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1365_1 ( .OUT(na1365_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na547_1), .IN5(1'b0), .IN6(na1265_1), .IN7(1'b0), .IN8(na1366_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1365_2 ( .OUT(na1365_1), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1365_1_i) );
// C_MX2b/D///      x156y64     80'h40_F800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_1 ( .OUT(na1366_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na547_1), .IN5(1'b0), .IN6(na1367_1), .IN7(1'b0), .IN8(na1857_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1366_2 ( .OUT(na1366_1), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1366_1_i) );
// C_MX2b/D///      x151y62     80'h40_F800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1367_1 ( .OUT(na1367_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na547_1), .IN5(1'b0), .IN6(na1286_1), .IN7(1'b0), .IN8(na1368_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1367_2 ( .OUT(na1367_1), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1367_1_i) );
// C_MX2b/D///      x152y62     80'h40_F800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1368_1 ( .OUT(na1368_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na547_1), .IN5(na1369_1), .IN6(1'b0), .IN7(na1297_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1368_2 ( .OUT(na1368_1), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1368_1_i) );
// C_MX2b/D///      x151y63     80'h40_F800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1369_1 ( .OUT(na1369_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na547_1), .IN5(na1150_2), .IN6(1'b0), .IN7(na1308_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1369_2 ( .OUT(na1369_1), .CLK(1'b0), .EN(na1395_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1369_1_i) );
// C_///AND/D      x147y59     80'h40_F800_80_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1370_4 ( .OUT(na1370_2_i), .IN1(~na1370_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1371_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1370_5 ( .OUT(na1370_2), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1370_2_i) );
// C_MX4a////      x148y60     80'h00_0018_00_0040_0CD9_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1371_1 ( .OUT(na1371_1), .IN1(~na4345_2), .IN2(1'b0), .IN3(1'b1), .IN4(~na1386_2), .IN5(na3235_2), .IN6(1'b1), .IN7(na1372_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y59     80'h00_0018_00_0000_0888_4282
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1372_1 ( .OUT(na1372_1), .IN1(na1377_1), .IN2(~na1383_1), .IN3(na1379_1), .IN4(na1375_1), .IN5(na1377_2), .IN6(~na1383_2),
                      .IN7(~na1379_2), .IN8(na1376_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y60     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1375_1 ( .OUT(na1375_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1370_2), .IN6(~na1378_1), .IN7(~na1380_1),
                      .IN8(~na1382_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x150y62     80'h40_F800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1376_1 ( .OUT(na1376_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1902_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1371_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1376_2 ( .OUT(na1376_1), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1376_1_i) );
// C_AND/D//AND/D      x151y61     80'h40_F800_80_0000_0C88_3A3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1377_1 ( .OUT(na1377_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1902_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1371_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1377_2 ( .OUT(na1377_1), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1377_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1377_4 ( .OUT(na1377_2_i), .IN1(na1906_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1371_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1377_5 ( .OUT(na1377_2), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1377_2_i) );
// C_AND/D///      x149y62     80'h40_F800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1378_1 ( .OUT(na1378_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1904_1), .IN7(1'b1), .IN8(~na1371_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1378_2 ( .OUT(na1378_1), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1378_1_i) );
// C_AND/D//AND/D      x150y65     80'h40_F800_80_0000_0C88_3C3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1379_1 ( .OUT(na1379_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1904_2), .IN7(1'b1), .IN8(~na1371_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1379_2 ( .OUT(na1379_1), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1379_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1379_4 ( .OUT(na1379_2_i), .IN1(na1910_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1371_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1379_5 ( .OUT(na1379_2), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1379_2_i) );
// C_AND/D///      x150y63     80'h40_F800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1380_1 ( .OUT(na1380_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1906_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1371_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1380_2 ( .OUT(na1380_1), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1380_1_i) );
// C_///AND/D      x150y62     80'h40_F800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1382_4 ( .OUT(na1382_2_i), .IN1(1'b1), .IN2(na1908_1), .IN3(1'b1), .IN4(~na1371_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1382_5 ( .OUT(na1382_2), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1382_2_i) );
// C_AND/D//AND/D      x149y64     80'h40_F800_80_0000_0C88_3C3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1383_1 ( .OUT(na1383_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1908_2), .IN7(1'b1), .IN8(~na1371_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1383_2 ( .OUT(na1383_1), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1383_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1383_4 ( .OUT(na1383_2_i), .IN1(na1910_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1371_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1383_5 ( .OUT(na1383_2), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1383_2_i) );
// C_///XOR/D      x154y60     80'h40_E800_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1386_4 ( .OUT(na1386_2_i), .IN1(na3235_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1386_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1386_5 ( .OUT(na1386_2), .CLK(1'b0), .EN(na1391_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1386_2_i) );
// C_AND////D      x102y67     80'h40_E418_00_0000_0888_F53C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1), .IN1(1'b1), .IN2(na1337_1), .IN3(1'b1), .IN4(~na549_1), .IN5(~na539_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1387_5 ( .OUT(na1387_2), .CLK(1'b0), .EN(~na1470_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1387_1) );
// C_///AND/      x95y81     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1388_4 ( .OUT(na1388_2), .IN1(~na3_1), .IN2(~na5_2), .IN3(na1390_2), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y84     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1389_1 ( .OUT(na1389_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6_1), .IN6(~na5_1), .IN7(na1387_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y79     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1390_4 ( .OUT(na1390_2), .IN1(~na3_2), .IN2(1'b1), .IN3(na2_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x152y60     80'h00_0018_00_0040_0A50_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1391_1 ( .OUT(na1391_1), .IN1(na1392_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na547_1), .IN5(na548_2), .IN6(1'b0), .IN7(na1372_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y61     80'h00_0060_00_0000_0C08_FFC1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1392_4 ( .OUT(na1392_2), .IN1(~na3235_2), .IN2(~na1393_1), .IN3(1'b1), .IN4(na1386_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x151y64     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1393_1 ( .OUT(na1393_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4329_2), .IN6(na1216_2), .IN7(na1217_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y73     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1394_1 ( .OUT(na1394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1339_1), .IN6(na1361_1), .IN7(~na3196_2),
                      .IN8(na3289_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y62     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1395_1 ( .OUT(na1395_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1396_1), .IN7(~na3701_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x151y60     80'h00_0018_00_0000_0888_BFA5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1396_1 ( .OUT(na1396_1), .IN1(~na3235_2), .IN2(1'b0), .IN3(na3289_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na1372_1),
                      .IN8(~na1386_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x80y60     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1397_4 ( .OUT(na1397_2), .IN1(na4084_2), .IN2(na1398_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x83y60     80'h00_0018_00_0040_0CCB_5300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1398_1 ( .OUT(na1398_1), .IN1(na3223_1), .IN2(na1348_1), .IN3(1'b1), .IN4(~na4368_2), .IN5(1'b1), .IN6(~na1361_1), .IN7(~na3196_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x107y72     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1399_4 ( .OUT(na1399_2), .IN1(1'b1), .IN2(na1402_1), .IN3(na1401_2), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y78     80'h00_0018_00_0000_0C88_A2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1400_1 ( .OUT(na1400_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6_1), .IN6(~na5_1), .IN7(na1387_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x86y79     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1401_4 ( .OUT(na1401_2), .IN1(na3_2), .IN2(1'b1), .IN3(na2_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y80     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1402_1 ( .OUT(na1402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3_1), .IN6(na5_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x107y73     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1403_4 ( .OUT(na1403_2), .IN1(1'b1), .IN2(na1402_1), .IN3(na1390_2), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y74     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1404_1 ( .OUT(na1404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1402_1), .IN7(na1405_1), .IN8(na1400_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y77     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1405_1 ( .OUT(na1405_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3_2), .IN6(1'b1), .IN7(~na2_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x102y71     80'h00_0060_00_0000_0C08_FF44
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1406_4 ( .OUT(na1406_2), .IN1(~na3_2), .IN2(na1402_1), .IN3(~na2_1), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y76     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1407_4 ( .OUT(na1407_2), .IN1(1'b1), .IN2(na1408_1), .IN3(na1401_2), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y82     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1408_1 ( .OUT(na1408_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_1), .IN6(na5_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y76     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1409_1 ( .OUT(na1409_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1408_1), .IN7(na1390_2), .IN8(na1400_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x102y74     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1410_4 ( .OUT(na1410_2), .IN1(1'b1), .IN2(na1408_1), .IN3(na1405_1), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y74     80'h00_0018_00_0000_0C88_44FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_1 ( .OUT(na1411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_2), .IN6(na1408_1), .IN7(~na2_1), .IN8(na1400_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y76     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1412_1 ( .OUT(na1412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1413_2), .IN7(na1401_2), .IN8(na1400_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y78     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1413_4 ( .OUT(na1413_2), .IN1(na3_1), .IN2(~na5_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x105y76     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1414_4 ( .OUT(na1414_2), .IN1(1'b1), .IN2(na1413_2), .IN3(na1390_2), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x103y74     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1415_4 ( .OUT(na1415_2), .IN1(1'b1), .IN2(na1413_2), .IN3(na1405_1), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y71     80'h00_0060_00_0000_0C08_FF44
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1416_4 ( .OUT(na1416_2), .IN1(~na3_2), .IN2(na1413_2), .IN3(~na2_1), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y77     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1417_1 ( .OUT(na1417_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_1), .IN6(~na5_2), .IN7(na1401_2), .IN8(na1400_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y87     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1418_1 ( .OUT(na1418_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1408_1), .IN7(na1401_2), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y80     80'h00_0018_00_0000_0C88_A4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1419_1 ( .OUT(na1419_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6_1), .IN6(na5_1), .IN7(na1387_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y73     80'h00_0018_00_0000_0C88_44FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1420_1 ( .OUT(na1420_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_2), .IN6(na1402_1), .IN7(~na2_1), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x86y72     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1421_4 ( .OUT(na1421_2), .IN1(1'b1), .IN2(na1402_1), .IN3(na1405_1), .IN4(na1419_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y77     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1422_1 ( .OUT(na1422_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1402_1), .IN7(na1390_2), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y70     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1423_1 ( .OUT(na1423_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4347_2), .IN8(na543_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y74     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1424_1 ( .OUT(na1424_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_1), .IN6(~na5_2), .IN7(na1405_1), .IN8(na1400_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x102y76     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1425_4 ( .OUT(na1425_2), .IN1(~na3_1), .IN2(~na5_2), .IN3(na1390_2), .IN4(na1400_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x103y83     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1426_4 ( .OUT(na1426_2), .IN1(1'b1), .IN2(na1408_1), .IN3(na1390_2), .IN4(na1419_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y79     80'h00_0018_00_0000_0C88_44FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1427_1 ( .OUT(na1427_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_2), .IN6(na1413_2), .IN7(~na2_1), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y77     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1428_4 ( .OUT(na1428_2), .IN1(1'b1), .IN2(na1413_2), .IN3(na1405_1), .IN4(na1419_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y84     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1429_1 ( .OUT(na1429_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1413_2), .IN7(na1390_2), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y80     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1430_4 ( .OUT(na1430_2), .IN1(1'b1), .IN2(na1413_2), .IN3(na1401_2), .IN4(na1419_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y75     80'h00_0060_00_0000_0C08_FF44
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1431_4 ( .OUT(na1431_2), .IN1(~na3_2), .IN2(na1408_1), .IN3(~na2_1), .IN4(na1419_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y78     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1432_1 ( .OUT(na1432_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1408_1), .IN7(na1405_1), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y86     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1433_1 ( .OUT(na1433_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_1), .IN6(~na5_2), .IN7(na1401_2), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y79     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1434_4 ( .OUT(na1434_2), .IN1(1'b1), .IN2(na1402_1), .IN3(na1405_1), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x105y81     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1435_4 ( .OUT(na1435_2), .IN1(1'b1), .IN2(na1402_1), .IN3(na1390_2), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y86     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1436_1 ( .OUT(na1436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1402_1), .IN7(na1401_2), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y73     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1437_4 ( .OUT(na1437_2), .IN1(1'b1), .IN2(1'b1), .IN3(na4348_2), .IN4(na543_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y77     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1438_4 ( .OUT(na1438_2), .IN1(~na3_1), .IN2(~na5_2), .IN3(na1405_1), .IN4(na1419_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y83     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1439_1 ( .OUT(na1439_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_1), .IN6(~na5_2), .IN7(na1390_2), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y74     80'h00_0060_00_0000_0C08_FF44
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1440_4 ( .OUT(na1440_2), .IN1(~na3_2), .IN2(na1402_1), .IN3(~na2_1), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x103y80     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1441_4 ( .OUT(na1441_2), .IN1(1'b1), .IN2(na1413_2), .IN3(na1390_2), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y86     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1442_1 ( .OUT(na1442_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1413_2), .IN7(na1401_2), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y80     80'h00_0018_00_0000_0C88_44FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1443_1 ( .OUT(na1443_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_2), .IN6(na1408_1), .IN7(~na2_1), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y81     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1444_1 ( .OUT(na1444_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1408_1), .IN7(na1405_1), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x102y81     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1445_4 ( .OUT(na1445_2), .IN1(1'b1), .IN2(na1408_1), .IN3(na1390_2), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y87     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1446_1 ( .OUT(na1446_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1408_1), .IN7(na1401_2), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y80     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1447_1 ( .OUT(na1447_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1413_2), .IN7(na1405_1), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x89y64     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1448_4 ( .OUT(na1448_2), .IN1(na1339_1), .IN2(~na1361_1), .IN3(~na3196_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y62     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1449_1 ( .OUT(na1449_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1361_1), .IN7(na3196_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y77     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1450_4 ( .OUT(na1450_2), .IN1(~na552_2), .IN2(1'b1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x140y70     80'h00_0078_00_0000_0C88_F2F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3871_2), .IN6(~na1333_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1451_4 ( .OUT(na1451_2), .IN1(na16_2), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y79     80'h00_0018_00_0040_0C66_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1452_1 ( .OUT(na1452_1), .IN1(1'b0), .IN2(~na1333_2), .IN3(~na4176_2), .IN4(1'b0), .IN5(na21_1), .IN6(1'b1), .IN7(na1142_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x131y76     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1453_1 ( .OUT(na1453_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1454_1), .IN6(1'b0), .IN7(na349_2), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y79     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1454_1 ( .OUT(na1454_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_1), .IN5(~na552_2), .IN6(1'b0), .IN7(~na1142_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x136y83     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1455_1 ( .OUT(na1455_1), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4088_2), .IN6(na1333_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x144y83     80'h00_0060_00_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1456_4 ( .OUT(na1456_2), .IN1(~na21_1), .IN2(na1333_1), .IN3(na4089_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x140y83     80'h00_0018_00_0040_0C1D_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1458_1 ( .OUT(na1458_1), .IN1(~na552_2), .IN2(1'b0), .IN3(na1142_1), .IN4(na4091_1), .IN5(1'b1), .IN6(~na1333_2), .IN7(na4171_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x139y85     80'h00_0018_00_0040_0C06_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1459_1 ( .OUT(na1459_1), .IN1(1'b0), .IN2(na1333_1), .IN3(na1142_1), .IN4(1'b0), .IN5(~na4174_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x137y80     80'h00_0060_00_0000_0C08_FFCD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1460_4 ( .OUT(na1460_2), .IN1(~na21_1), .IN2(na1333_1), .IN3(1'b0), .IN4(na1461_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x128y68     80'h00_0018_00_0040_0C0C_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1461_1 ( .OUT(na1461_1), .IN1(1'b0), .IN2(1'b0), .IN3(na4093_1), .IN4(na1332_1), .IN5(~na1331_1), .IN6(1'b1), .IN7(~na4365_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x125y79     80'h00_0018_00_0040_0C1D_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1462_1 ( .OUT(na1462_1), .IN1(~na552_2), .IN2(1'b0), .IN3(na1142_1), .IN4(na4091_1), .IN5(1'b1), .IN6(~na1333_2), .IN7(1'b1),
                      .IN8(~na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x127y74     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1463_4 ( .OUT(na1463_2), .IN1(~na21_1), .IN2(~na4315_2), .IN3(1'b0), .IN4(~na4352_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y94     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1464_1 ( .OUT(na1464_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3871_2), .IN6(na1333_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x141y90     80'h00_0018_00_0000_0C88_D3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1465_1 ( .OUT(na1465_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1464_1), .IN7(~na1142_1), .IN8(na25_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x138y81     80'h00_0018_00_0000_0888_FE35
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1466_1 ( .OUT(na1466_1), .IN1(~na21_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na1451_1), .IN5(na552_2), .IN6(na4349_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y82     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1467_4 ( .OUT(na1467_2), .IN1(~na542_2), .IN2(~na1337_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x153y65     80'h00_0018_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1468_1 ( .OUT(na1468_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na539_1), .IN6(na545_2), .IN7(1'b0), .IN8(na549_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y80     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1469_1 ( .OUT(na1469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na25_2), .IN5(na4351_2), .IN6(1'b0), .IN7(na1142_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x140y63     80'h00_0060_00_0000_0C08_FFD3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1470_4 ( .OUT(na1470_2), .IN1(1'b0), .IN2(~na1399_2), .IN3(~na4202_2), .IN4(na549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y72     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1471_4 ( .OUT(na1471_2), .IN1(~na552_2), .IN2(1'b1), .IN3(~na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x133y84     80'h00_0018_00_0040_0C06_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1472_1 ( .OUT(na1472_1), .IN1(1'b0), .IN2(na1333_1), .IN3(na1142_1), .IN4(1'b0), .IN5(~na21_1), .IN6(1'b1), .IN7(1'b1), .IN8(na25_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x105y80     80'h00_0018_00_0000_0888_DF35
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1473_1 ( .OUT(na1473_1), .IN1(~na21_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na1471_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na4431_2),
                      .IN8(na1451_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y82     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1474_1 ( .OUT(na1474_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1402_1), .IN7(na1401_2), .IN8(na1419_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x103y82     80'h00_0018_00_0000_0888_DF5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1475_1 ( .OUT(na1475_1), .IN1(na552_2), .IN2(na4103_2), .IN3(~na4173_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(~na4431_2),
                      .IN8(na1451_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y76     80'h00_0060_00_0000_0C08_FF44
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1477_4 ( .OUT(na1477_2), .IN1(~na3_2), .IN2(na1413_2), .IN3(~na2_1), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y85     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1478_1 ( .OUT(na1478_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_1), .IN6(~na5_2), .IN7(na1401_2), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y78     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1479_4 ( .OUT(na1479_2), .IN1(1'b1), .IN2(1'b1), .IN3(na4346_2), .IN4(na543_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y80     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1480_4 ( .OUT(na1480_2), .IN1(~na3_1), .IN2(~na5_2), .IN3(na1405_1), .IN4(na1389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x143y61     80'h00_0018_00_0040_0C05_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1481_1 ( .OUT(na1481_1), .IN1(na4105_2), .IN2(1'b0), .IN3(na4104_1), .IN4(1'b0), .IN5(na3142_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na3144_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x107y100     80'hC0_EC18_00_0000_0666_AC3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1482_1 ( .OUT(na1482_1), .IN1(na1014_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na640_1), .IN5(1'b0), .IN6(na973_1), .IN7(na809_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1482_5 ( .OUT(na1482_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1482_1) );
// C_XOR////D      x109y99     80'hC0_EC18_00_0000_0666_59C0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1483_1 ( .OUT(na1483_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1022_2), .IN5(na1019_1), .IN6(~na641_1), .IN7(~na808_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1483_5 ( .OUT(na1483_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1483_1) );
// C_XOR////D      x117y101     80'hC0_EC18_00_0000_0666_CC9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1484_1 ( .OUT(na1484_1), .IN1(na810_2), .IN2(1'b0), .IN3(~na1033_1), .IN4(na1031_1), .IN5(1'b0), .IN6(na973_1), .IN7(1'b0),
                      .IN8(na642_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1484_5 ( .OUT(na1484_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1484_1) );
// C_XOR////D      x104y97     80'hC0_EC18_00_0000_0666_069A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1486_1 ( .OUT(na1486_1), .IN1(na643_1), .IN2(1'b0), .IN3(na1033_1), .IN4(~na1036_1), .IN5(na811_1), .IN6(na973_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1486_5 ( .OUT(na1486_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1486_1) );
// C_XOR////D      x106y97     80'hC0_EC18_00_0000_0666_63CA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1488_1 ( .OUT(na1488_1), .IN1(na812_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1036_1), .IN5(1'b0), .IN6(~na1042_2), .IN7(na1033_1),
                      .IN8(na644_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1488_5 ( .OUT(na1488_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1488_1) );
// C_XOR////D      x91y95     80'hC0_EC18_00_0000_0666_6CC5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1490_1 ( .OUT(na1490_1), .IN1(~na1026_1), .IN2(1'b0), .IN3(1'b0), .IN4(na813_1), .IN5(1'b0), .IN6(na1046_1), .IN7(na1047_1),
                      .IN8(na645_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1490_5 ( .OUT(na1490_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1490_1) );
// C_XOR////D      x90y82     80'hC0_EC18_00_0000_0666_9090
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1492_1 ( .OUT(na1492_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1023_2), .IN4(~na646_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1047_1),
                      .IN8(~na814_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1492_5 ( .OUT(na1492_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1492_1) );
// C_XOR////D      x85y76     80'hC0_EC18_00_0000_0666_C063
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1493_1 ( .OUT(na1493_1), .IN1(1'b0), .IN2(~na647_1), .IN3(na1047_1), .IN4(na815_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1022_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1493_5 ( .OUT(na1493_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1493_1) );
// C_XOR////D      x88y81     80'hC0_EC18_00_0000_0666_A0C0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1494_1 ( .OUT(na1494_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na616_1), .IN5(1'b0), .IN6(1'b0), .IN7(na214_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1494_5 ( .OUT(na1494_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1494_1) );
// C_///XOR/D      x114y75     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1495_4 ( .OUT(na1495_2_i), .IN1(na264_1), .IN2(1'b0), .IN3(na617_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1495_5 ( .OUT(na1495_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1495_2_i) );
// C_XOR/D///      x116y85     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1496_1 ( .OUT(na1496_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na618_1), .IN6(1'b0), .IN7(1'b0), .IN8(na277_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1496_2 ( .OUT(na1496_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1496_1_i) );
// C_XOR/D///      x114y64     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1497_1 ( .OUT(na1497_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na619_1), .IN7(na287_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1497_2 ( .OUT(na1497_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1497_1_i) );
// C_XOR/D///      x93y64     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1498_1 ( .OUT(na1498_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na295_1), .IN8(na620_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1498_2 ( .OUT(na1498_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1498_1_i) );
// C_XOR////D      x84y68     80'hC0_EC18_00_0000_0666_09A0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1499_1 ( .OUT(na1499_1), .IN1(1'b0), .IN2(1'b0), .IN3(na301_2), .IN4(1'b0), .IN5(~na621_1), .IN6(na303_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1499_5 ( .OUT(na1499_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1499_1) );
// C_XOR////D      x86y59     80'hC0_EC18_00_0000_0666_60A0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1500_1 ( .OUT(na1500_1), .IN1(1'b0), .IN2(1'b0), .IN3(na622_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na301_2), .IN8(na310_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1500_5 ( .OUT(na1500_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1500_1) );
// C_///XOR/D      x109y60     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1501_4 ( .OUT(na1501_2_i), .IN1(na315_1), .IN2(na623_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1501_5 ( .OUT(na1501_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1501_2_i) );
// C_XOR////D      x87y84     80'hC0_EC18_00_0000_0666_0CCC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1502_1 ( .OUT(na1502_1), .IN1(1'b0), .IN2(na817_1), .IN3(1'b0), .IN4(na624_1), .IN5(1'b0), .IN6(na855_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1502_5 ( .OUT(na1502_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1502_1) );
// C_XOR/D///      x104y90     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1503_1 ( .OUT(na1503_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na625_1), .IN6(na862_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1503_2 ( .OUT(na1503_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1503_1_i) );
// C_XOR////D      x94y96     80'hC0_EC18_00_0000_0666_0C9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1504_1 ( .OUT(na1504_1), .IN1(na872_1), .IN2(1'b0), .IN3(~na874_1), .IN4(na626_1), .IN5(1'b0), .IN6(na873_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1504_5 ( .OUT(na1504_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1504_1) );
// C_///XOR/D      x112y70     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1505_4 ( .OUT(na1505_2_i), .IN1(na627_1), .IN2(na877_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1505_5 ( .OUT(na1505_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1505_2_i) );
// C_///XOR/D      x97y74     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1506_4 ( .OUT(na1506_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na628_1), .IN4(na883_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1506_5 ( .OUT(na1506_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1506_2_i) );
// C_XOR////D      x82y77     80'hC0_EC18_00_0000_0666_AC35
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1507_1 ( .OUT(na1507_1), .IN1(~na875_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na629_1), .IN5(1'b0), .IN6(na817_1), .IN7(na888_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1507_5 ( .OUT(na1507_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1507_1) );
// C_XOR////D      x82y66     80'hC0_EC18_00_0000_0666_6030
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1508_1 ( .OUT(na1508_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(~na630_1), .IN5(1'b0), .IN6(1'b0), .IN7(na888_1), .IN8(na864_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1508_5 ( .OUT(na1508_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1508_1) );
// C_XOR////D      x83y63     80'hC0_EC18_00_0000_0666_AA0C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1509_1 ( .OUT(na1509_1), .IN1(1'b0), .IN2(na631_1), .IN3(1'b0), .IN4(1'b0), .IN5(na893_2), .IN6(1'b0), .IN7(na888_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1509_5 ( .OUT(na1509_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1509_1) );
// C_///XOR/D      x138y97     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1510_4 ( .OUT(na1510_2_i), .IN1(na632_1), .IN2(1'b0), .IN3(1'b0), .IN4(na895_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1510_5 ( .OUT(na1510_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1510_2_i) );
// C_XOR/D///      x131y101     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1511_1 ( .OUT(na1511_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na633_1), .IN7(na4285_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1511_2 ( .OUT(na1511_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1511_1_i) );
// C_XOR////D      x133y102     80'hC0_EC18_00_0000_0666_AC5A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1512_1 ( .OUT(na1512_1), .IN1(na634_1), .IN2(1'b0), .IN3(~na952_1), .IN4(1'b0), .IN5(1'b0), .IN6(na950_1), .IN7(na951_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1512_5 ( .OUT(na1512_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1512_1) );
// C_XOR////D      x139y98     80'hC0_EC18_00_0000_0666_6035
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1513_1 ( .OUT(na1513_1), .IN1(~na957_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na635_1), .IN5(1'b0), .IN6(1'b0), .IN7(na952_1), .IN8(na956_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1513_5 ( .OUT(na1513_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1513_1) );
// C_XOR/D///      x144y93     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1514_1 ( .OUT(na1514_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na636_1), .IN7(na962_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1514_2 ( .OUT(na1514_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1514_1_i) );
// C_XOR/D///      x123y87     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1515_1 ( .OUT(na1515_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na965_1), .IN7(1'b0), .IN8(na637_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1515_2 ( .OUT(na1515_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1515_1_i) );
// C_XOR////D      x117y64     80'hC0_EC18_00_0000_0666_A00C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1516_1 ( .OUT(na1516_1), .IN1(1'b0), .IN2(na968_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na638_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1516_5 ( .OUT(na1516_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1516_1) );
// C_///XOR/D      x136y67     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1517_4 ( .OUT(na1517_2_i), .IN1(na970_1), .IN2(1'b0), .IN3(na639_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1517_5 ( .OUT(na1517_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1517_2_i) );
// C_///XOR/D      x83y78     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1518_4 ( .OUT(na1518_2_i), .IN1(na648_1), .IN2(1'b0), .IN3(na1494_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1518_5 ( .OUT(na1518_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1518_2_i) );
// C_///XOR/D      x119y84     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1519_4 ( .OUT(na1519_2_i), .IN1(na264_1), .IN2(1'b0), .IN3(na617_1), .IN4(na649_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1519_5 ( .OUT(na1519_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1519_2_i) );
// C_XOR/D///      x119y87     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1520_1 ( .OUT(na1520_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na618_1), .IN6(1'b0), .IN7(na650_1), .IN8(na277_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1520_2 ( .OUT(na1520_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1520_1_i) );
// C_///XOR/D      x115y62     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1521_4 ( .OUT(na1521_2_i), .IN1(na651_1), .IN2(na619_1), .IN3(na287_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1521_5 ( .OUT(na1521_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1521_2_i) );
// C_///XOR/D      x92y65     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1522_4 ( .OUT(na1522_2_i), .IN1(na652_1), .IN2(1'b0), .IN3(na295_1), .IN4(na620_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1522_5 ( .OUT(na1522_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1522_2_i) );
// C_///XOR/D      x83y65     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1523_4 ( .OUT(na1523_2_i), .IN1(na653_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1499_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1523_5 ( .OUT(na1523_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1523_2_i) );
// C_XOR/D///      x88y58     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1524_1 ( .OUT(na1524_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1500_1), .IN8(na654_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1524_2 ( .OUT(na1524_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1524_1_i) );
// C_///XOR/D      x104y63     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1525_4 ( .OUT(na1525_2_i), .IN1(na315_1), .IN2(na623_1), .IN3(1'b0), .IN4(na655_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1525_5 ( .OUT(na1525_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1525_2_i) );
// C_XOR/D///      x89y84     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1526_1 ( .OUT(na1526_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1502_1), .IN7(1'b0), .IN8(na656_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1526_2 ( .OUT(na1526_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1526_1_i) );
// C_XOR/D///      x101y87     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1527_1 ( .OUT(na1527_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na625_1), .IN6(na862_1), .IN7(1'b0), .IN8(na657_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1527_2 ( .OUT(na1527_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1527_1_i) );
// C_XOR/D///      x95y95     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1528_1 ( .OUT(na1528_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na658_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1504_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1528_2 ( .OUT(na1528_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1528_1_i) );
// C_XOR////D      x92y81     80'hC0_EC18_00_0000_0666_CA09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1529_1 ( .OUT(na1529_1), .IN1(na627_1), .IN2(~na659_1), .IN3(1'b0), .IN4(1'b0), .IN5(na872_1), .IN6(1'b0), .IN7(1'b0), .IN8(na878_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1529_5 ( .OUT(na1529_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1529_1) );
// C_XOR////D      x87y82     80'hC0_EC18_00_0000_0666_CC53
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1530_1 ( .OUT(na1530_1), .IN1(1'b0), .IN2(~na660_1), .IN3(~na628_1), .IN4(1'b0), .IN5(1'b0), .IN6(na884_2), .IN7(1'b0), .IN8(na878_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1530_5 ( .OUT(na1530_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1530_1) );
// C_///XOR/D      x81y70     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1531_4 ( .OUT(na1531_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1507_1), .IN4(na661_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1531_5 ( .OUT(na1531_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1531_2_i) );
// C_///XOR/D      x85y65     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1532_4 ( .OUT(na1532_2_i), .IN1(na662_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1508_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1532_5 ( .OUT(na1532_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1532_2_i) );
// C_///XOR/D      x90y60     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1533_4 ( .OUT(na1533_2_i), .IN1(na1509_1), .IN2(1'b0), .IN3(na663_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1533_5 ( .OUT(na1533_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1533_2_i) );
// C_///XOR/D      x139y100     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1534_4 ( .OUT(na1534_2_i), .IN1(na632_1), .IN2(na664_1), .IN3(1'b0), .IN4(na895_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1534_5 ( .OUT(na1534_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1534_2_i) );
// C_///XOR/D      x134y99     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1535_4 ( .OUT(na1535_2_i), .IN1(na665_1), .IN2(na633_1), .IN3(na4285_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1535_5 ( .OUT(na1535_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1535_2_i) );
// C_XOR/D///      x127y103     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1536_1 ( .OUT(na1536_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1512_1), .IN7(1'b0), .IN8(na666_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1536_2 ( .OUT(na1536_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1536_1_i) );
// C_XOR/D///      x139y95     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1537_1 ( .OUT(na1537_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1513_1), .IN7(na667_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1537_2 ( .OUT(na1537_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1537_1_i) );
// C_XOR////D      x137y94     80'hC0_EC18_00_0000_0666_AA5C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1538_1 ( .OUT(na1538_1), .IN1(1'b0), .IN2(na636_1), .IN3(~na668_1), .IN4(1'b0), .IN5(na963_1), .IN6(1'b0), .IN7(na952_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1538_5 ( .OUT(na1538_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1538_1) );
// C_XOR////D      x119y89     80'hC0_EC18_00_0000_0666_A33A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1539_1 ( .OUT(na1539_1), .IN1(na963_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na637_1), .IN5(1'b0), .IN6(~na669_1), .IN7(na966_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1539_5 ( .OUT(na1539_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1539_1) );
// C_XOR/D///      x111y63     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1540_1 ( .OUT(na1540_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na670_1), .IN6(na1516_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1540_2 ( .OUT(na1540_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1540_1_i) );
// C_XOR////D      x131y79     80'hC0_EC18_00_0000_0666_AA53
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1541_1 ( .OUT(na1541_1), .IN1(1'b0), .IN2(~na671_1), .IN3(~na639_1), .IN4(1'b0), .IN5(na963_1), .IN6(1'b0), .IN7(na951_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1541_5 ( .OUT(na1541_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1541_1) );
// C_///XOR/D      x111y98     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1542_4 ( .OUT(na1542_2_i), .IN1(1'b0), .IN2(na1482_1), .IN3(1'b0), .IN4(na672_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1542_5 ( .OUT(na1542_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1542_2_i) );
// C_///XOR/D      x113y102     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1543_4 ( .OUT(na1543_2_i), .IN1(na1483_1), .IN2(na673_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1543_5 ( .OUT(na1543_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1543_2_i) );
// C_///XOR/D      x119y102     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1544_4 ( .OUT(na1544_2_i), .IN1(na1484_1), .IN2(na674_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1544_5 ( .OUT(na1544_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1544_2_i) );
// C_XOR/D///      x99y96     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1545_1 ( .OUT(na1545_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na675_1), .IN7(na1486_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1545_2 ( .OUT(na1545_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1545_1_i) );
// C_///XOR/D      x93y93     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1546_4 ( .OUT(na1546_2_i), .IN1(1'b0), .IN2(na676_1), .IN3(na1488_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1546_5 ( .OUT(na1546_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1546_2_i) );
// C_XOR/D///      x94y91     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1547_1 ( .OUT(na1547_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1490_1), .IN6(1'b0), .IN7(1'b0), .IN8(na677_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1547_2 ( .OUT(na1547_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1547_1_i) );
// C_XOR/D///      x88y74     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1548_1 ( .OUT(na1548_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na678_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1492_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1548_2 ( .OUT(na1548_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1548_1_i) );
// C_XOR/D///      x87y70     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1549_1 ( .OUT(na1549_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na679_1), .IN6(na1493_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1549_2 ( .OUT(na1549_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1549_1_i) );
// C_XOR/D///      x91y85     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1550_1 ( .OUT(na1550_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na648_1), .IN6(1'b0), .IN7(na1494_1), .IN8(na680_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1550_2 ( .OUT(na1550_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1550_1_i) );
// C_XOR/D///      x114y79     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1551_1 ( .OUT(na1551_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na264_1), .IN6(na681_1), .IN7(~na617_1),
                      .IN8(~na649_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1551_2 ( .OUT(na1551_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1551_1_i) );
// C_///XOR/D      x117y88     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1552_4 ( .OUT(na1552_2_i), .IN1(~na618_1), .IN2(na682_1), .IN3(~na650_1), .IN4(na277_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1552_5 ( .OUT(na1552_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1552_2_i) );
// C_XOR/D///      x112y63     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1553_1 ( .OUT(na1553_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na651_1), .IN6(~na619_1), .IN7(na287_1),
                      .IN8(na683_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1553_2 ( .OUT(na1553_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1553_1_i) );
// C_XOR/D///      x99y67     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1554_1 ( .OUT(na1554_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na652_1), .IN6(na684_1), .IN7(na295_1),
                      .IN8(~na620_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1554_2 ( .OUT(na1554_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1554_1_i) );
// C_///XOR/D      x85y66     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1555_4 ( .OUT(na1555_2_i), .IN1(na653_1), .IN2(1'b0), .IN3(na685_1), .IN4(na1499_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1555_5 ( .OUT(na1555_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1555_2_i) );
// C_XOR/D///      x90y59     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1556_1 ( .OUT(na1556_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na686_1), .IN7(na1500_1), .IN8(na654_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1556_2 ( .OUT(na1556_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1556_1_i) );
// C_XOR/D///      x101y59     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1557_1 ( .OUT(na1557_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na315_1), .IN6(~na623_1), .IN7(na687_1),
                      .IN8(~na655_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1557_2 ( .OUT(na1557_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1557_1_i) );
// C_///XOR/D      x87y81     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1558_4 ( .OUT(na1558_2_i), .IN1(1'b0), .IN2(na1502_1), .IN3(na688_1), .IN4(na656_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1558_5 ( .OUT(na1558_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1558_2_i) );
// C_XOR/D///      x105y92     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1559_1 ( .OUT(na1559_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na625_1), .IN6(na862_1), .IN7(na689_1),
                      .IN8(~na657_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1559_2 ( .OUT(na1559_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1559_1_i) );
// C_XOR/D///      x97y96     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1560_1 ( .OUT(na1560_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na658_1), .IN6(1'b0), .IN7(na690_1), .IN8(na1504_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1560_2 ( .OUT(na1560_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1560_1_i) );
// C_///XOR/D      x87y72     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1561_4 ( .OUT(na1561_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1529_1), .IN4(na691_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1561_5 ( .OUT(na1561_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1561_2_i) );
// C_///XOR/D      x87y73     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1562_4 ( .OUT(na1562_2_i), .IN1(1'b0), .IN2(na1530_1), .IN3(na692_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1562_5 ( .OUT(na1562_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1562_2_i) );
// C_///XOR/D      x81y69     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1563_4 ( .OUT(na1563_2_i), .IN1(1'b0), .IN2(na693_1), .IN3(na1507_1), .IN4(na661_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1563_5 ( .OUT(na1563_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1563_2_i) );
// C_XOR/D///      x85y65     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1564_1 ( .OUT(na1564_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na662_1), .IN6(na694_1), .IN7(1'b0), .IN8(na1508_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1564_2 ( .OUT(na1564_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1564_1_i) );
// C_///XOR/D      x93y61     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1565_4 ( .OUT(na1565_2_i), .IN1(na1509_1), .IN2(na695_1), .IN3(na663_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1565_5 ( .OUT(na1565_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1565_2_i) );
// C_///XOR/D      x136y97     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1566_4 ( .OUT(na1566_2_i), .IN1(~na632_1), .IN2(~na664_1), .IN3(na696_1), .IN4(na895_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1566_5 ( .OUT(na1566_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1566_2_i) );
// C_XOR/D///      x131y103     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1567_1 ( .OUT(na1567_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na665_1), .IN6(~na633_1), .IN7(na4285_2),
                      .IN8(na697_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1567_2 ( .OUT(na1567_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1567_1_i) );
// C_XOR/D///      x132y101     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1568_1 ( .OUT(na1568_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1512_1), .IN7(na698_1), .IN8(na666_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1568_2 ( .OUT(na1568_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1568_1_i) );
// C_///XOR/D      x135y96     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1569_4 ( .OUT(na1569_2_i), .IN1(1'b0), .IN2(na1513_1), .IN3(na667_1), .IN4(na699_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1569_5 ( .OUT(na1569_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1569_2_i) );
// C_///XOR/D      x131y87     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1570_4 ( .OUT(na1570_2_i), .IN1(1'b0), .IN2(na1538_1), .IN3(na700_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1570_5 ( .OUT(na1570_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1570_2_i) );
// C_XOR/D///      x113y94     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1571_1 ( .OUT(na1571_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1539_1), .IN6(1'b0), .IN7(na701_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1571_2 ( .OUT(na1571_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1571_1_i) );
// C_///XOR/D      x115y64     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1572_4 ( .OUT(na1572_2_i), .IN1(na670_1), .IN2(na702_1), .IN3(na4356_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1572_5 ( .OUT(na1572_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1572_2_i) );
// C_XOR/D///      x125y71     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1573_1 ( .OUT(na1573_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1541_1), .IN6(1'b0), .IN7(na703_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1573_2 ( .OUT(na1573_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1573_1_i) );
// C_XOR/D///      x113y97     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1574_1 ( .OUT(na1574_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1482_1), .IN7(na704_1), .IN8(na672_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1574_2 ( .OUT(na1574_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1574_1_i) );
// C_///XOR/D      x116y99     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1575_4 ( .OUT(na1575_2_i), .IN1(na1483_1), .IN2(na673_1), .IN3(1'b0), .IN4(na705_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1575_5 ( .OUT(na1575_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1575_2_i) );
// C_XOR/D///      x121y101     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1576_1 ( .OUT(na1576_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1484_1), .IN6(na674_1), .IN7(1'b0), .IN8(na706_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1576_2 ( .OUT(na1576_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1576_1_i) );
// C_///XOR/D      x97y93     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1577_4 ( .OUT(na1577_2_i), .IN1(1'b0), .IN2(na675_1), .IN3(na1486_1), .IN4(na707_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1577_5 ( .OUT(na1577_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1577_2_i) );
// C_XOR/D///      x97y93     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1578_1 ( .OUT(na1578_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na676_1), .IN7(na1488_1), .IN8(na708_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1578_2 ( .OUT(na1578_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1578_1_i) );
// C_///XOR/D      x87y85     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1579_4 ( .OUT(na1579_2_i), .IN1(na1490_1), .IN2(na709_1), .IN3(1'b0), .IN4(na677_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1579_5 ( .OUT(na1579_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1579_2_i) );
// C_XOR/D///      x87y72     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1580_1 ( .OUT(na1580_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na678_1), .IN6(na710_1), .IN7(1'b0), .IN8(na1492_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1580_2 ( .OUT(na1580_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1580_1_i) );
// C_///XOR/D      x87y67     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1581_4 ( .OUT(na1581_2_i), .IN1(na679_1), .IN2(na1493_1), .IN3(1'b0), .IN4(na711_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1581_5 ( .OUT(na1581_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1581_2_i) );
// C_///XOR/D      x89y84     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1582_4 ( .OUT(na1582_2_i), .IN1(~na648_1), .IN2(na551_1), .IN3(na1494_1), .IN4(~na680_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1582_5 ( .OUT(na1582_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1582_2_i) );
// C_XOR/D///      x115y81     80'hC0_EC00_00_0000_0666_3A56
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1583_1 ( .OUT(na1583_1_i), .IN1(na553_1), .IN2(na681_1), .IN3(~na617_1), .IN4(1'b0), .IN5(na264_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(~na649_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1583_2 ( .OUT(na1583_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1583_1_i) );
// C_XOR/D///      x114y88     80'hC0_EC00_00_0000_0666_CC59
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1584_1 ( .OUT(na1584_1_i), .IN1(~na618_1), .IN2(na682_1), .IN3(~na650_1), .IN4(1'b0), .IN5(1'b0), .IN6(na554_1), .IN7(1'b0),
                      .IN8(na277_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1584_2 ( .OUT(na1584_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1584_1_i) );
// C_XOR/D///      x107y65     80'hC0_EC00_00_0000_0666_AAC6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1585_1 ( .OUT(na1585_1_i), .IN1(~na651_1), .IN2(~na619_1), .IN3(1'b0), .IN4(na683_1), .IN5(na555_1), .IN6(1'b0), .IN7(na287_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1585_2 ( .OUT(na1585_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1585_1_i) );
// C_XOR/D///      x95y69     80'hC0_EC00_00_0000_0666_0A99
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1586_1 ( .OUT(na1586_1_i), .IN1(~na652_1), .IN2(na684_1), .IN3(na295_1), .IN4(~na620_1), .IN5(na556_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1586_2 ( .OUT(na1586_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1586_1_i) );
// C_///XOR/D      x83y69     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1587_4 ( .OUT(na1587_2_i), .IN1(~na653_1), .IN2(na557_1), .IN3(~na685_1), .IN4(na1499_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1587_5 ( .OUT(na1587_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1587_2_i) );
// C_///XOR/D      x97y61     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1588_4 ( .OUT(na1588_2_i), .IN1(na558_1), .IN2(~na686_1), .IN3(na1500_1), .IN4(~na654_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1588_5 ( .OUT(na1588_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1588_2_i) );
// C_XOR/D///      x102y63     80'hC0_EC00_00_0000_0666_AA93
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1589_1 ( .OUT(na1589_1_i), .IN1(1'b0), .IN2(~na623_1), .IN3(na687_1), .IN4(~na655_1), .IN5(na315_1), .IN6(1'b0), .IN7(na559_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1589_2 ( .OUT(na1589_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1589_1_i) );
// C_///XOR/D      x83y82     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1590_4 ( .OUT(na1590_2_i), .IN1(na560_1), .IN2(na1502_1), .IN3(~na688_1), .IN4(~na656_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1590_5 ( .OUT(na1590_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1590_2_i) );
// C_XOR/D///      x105y91     80'hC0_EC00_00_0000_0666_36A5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1591_1 ( .OUT(na1591_1_i), .IN1(~na625_1), .IN2(1'b0), .IN3(na689_1), .IN4(1'b0), .IN5(na561_1), .IN6(na862_1), .IN7(1'b0),
                      .IN8(~na657_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1591_2 ( .OUT(na1591_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1591_1_i) );
// C_XOR/D///      x97y94     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1592_1 ( .OUT(na1592_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na658_1), .IN6(na562_1), .IN7(~na690_1),
                      .IN8(na1504_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1592_2 ( .OUT(na1592_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1592_1_i) );
// C_XOR/D///      x97y79     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1593_1 ( .OUT(na1593_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na563_1), .IN6(1'b0), .IN7(na1529_1), .IN8(na691_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1593_2 ( .OUT(na1593_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1593_1_i) );
// C_XOR/D///      x88y80     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1594_1 ( .OUT(na1594_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na564_1), .IN6(na1530_1), .IN7(na692_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1594_2 ( .OUT(na1594_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1594_1_i) );
// C_///XOR/D      x83y71     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1595_4 ( .OUT(na1595_2_i), .IN1(na565_1), .IN2(~na693_1), .IN3(na1507_1), .IN4(~na661_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1595_5 ( .OUT(na1595_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1595_2_i) );
// C_XOR/D///      x86y65     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1596_1 ( .OUT(na1596_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na662_1), .IN6(~na694_1), .IN7(na566_1),
                      .IN8(na1508_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1596_2 ( .OUT(na1596_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1596_1_i) );
// C_///XOR/D      x93y64     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1597_4 ( .OUT(na1597_2_i), .IN1(na1509_1), .IN2(~na695_1), .IN3(~na663_1), .IN4(na567_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1597_5 ( .OUT(na1597_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1597_2_i) );
// C_XOR/D///      x131y98     80'hC0_EC00_00_0000_0666_CAA6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1598_1 ( .OUT(na1598_1_i), .IN1(~na632_1), .IN2(~na664_1), .IN3(na696_1), .IN4(1'b0), .IN5(na568_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na895_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1598_2 ( .OUT(na1598_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1598_1_i) );
// C_XOR/D///      x127y100     80'hC0_EC00_00_0000_0666_AAC6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_1 ( .OUT(na1599_1_i), .IN1(~na665_1), .IN2(~na633_1), .IN3(1'b0), .IN4(na697_1), .IN5(na569_1), .IN6(1'b0), .IN7(na4285_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1599_2 ( .OUT(na1599_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1599_1_i) );
// C_XOR/D///      x125y101     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1600_1 ( .OUT(na1600_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na570_1), .IN6(na1512_1), .IN7(~na698_1),
                      .IN8(~na666_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1600_2 ( .OUT(na1600_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1600_1_i) );
// C_///XOR/D      x136y95     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1601_4 ( .OUT(na1601_2_i), .IN1(na571_1), .IN2(na1513_1), .IN3(~na667_1), .IN4(~na699_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1601_5 ( .OUT(na1601_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1601_2_i) );
// C_///XOR/D      x123y89     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1602_4 ( .OUT(na1602_2_i), .IN1(na572_1), .IN2(na1538_1), .IN3(na700_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1602_5 ( .OUT(na1602_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1602_2_i) );
// C_///XOR/D      x113y90     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1603_4 ( .OUT(na1603_2_i), .IN1(na1539_1), .IN2(na573_1), .IN3(na701_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1603_5 ( .OUT(na1603_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1603_2_i) );
// C_///XOR/D      x112y63     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1604_4 ( .OUT(na1604_2_i), .IN1(~na670_1), .IN2(~na702_1), .IN3(na4356_2), .IN4(na574_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1604_5 ( .OUT(na1604_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1604_2_i) );
// C_XOR/D///      x125y72     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1605_1 ( .OUT(na1605_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1541_1), .IN6(1'b0), .IN7(na703_1), .IN8(na4212_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1605_2 ( .OUT(na1605_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1605_1_i) );
// C_///XOR/D      x103y95     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1606_4 ( .OUT(na1606_2_i), .IN1(na576_1), .IN2(na1482_1), .IN3(~na704_1), .IN4(~na672_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1606_5 ( .OUT(na1606_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1606_2_i) );
// C_XOR/D///      x116y99     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1607_1 ( .OUT(na1607_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1483_1), .IN6(~na673_1), .IN7(na577_1),
                      .IN8(~na705_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1607_2 ( .OUT(na1607_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1607_1_i) );
// C_///XOR/D      x118y100     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1608_4 ( .OUT(na1608_2_i), .IN1(na1484_1), .IN2(~na674_1), .IN3(na578_1), .IN4(~na706_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1608_5 ( .OUT(na1608_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1608_2_i) );
// C_XOR/D///      x101y91     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1609_1 ( .OUT(na1609_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na579_1), .IN6(~na675_1), .IN7(na1486_1),
                      .IN8(~na707_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1609_2 ( .OUT(na1609_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1609_1_i) );
// C_///XOR/D      x97y92     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1610_4 ( .OUT(na1610_2_i), .IN1(na580_1), .IN2(~na676_1), .IN3(na1488_1), .IN4(~na708_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1610_5 ( .OUT(na1610_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1610_2_i) );
// C_///XOR/D      x91y87     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1611_4 ( .OUT(na1611_2_i), .IN1(na1490_1), .IN2(~na709_1), .IN3(na581_1), .IN4(~na677_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1611_5 ( .OUT(na1611_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1611_2_i) );
// C_XOR/D///      x91y74     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1612_1 ( .OUT(na1612_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na678_1), .IN6(~na710_1), .IN7(na582_1),
                      .IN8(na1492_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1612_2 ( .OUT(na1612_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1612_1_i) );
// C_///XOR/D      x89y69     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1613_4 ( .OUT(na1613_2_i), .IN1(~na679_1), .IN2(na1493_1), .IN3(na583_1), .IN4(~na711_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1613_5 ( .OUT(na1613_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1613_2_i) );
// C_XOR////D      x92y85     80'hC0_EC18_00_0000_0666_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1614_1 ( .OUT(na1614_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na712_1), .IN7(na214_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1614_5 ( .OUT(na1614_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1614_1) );
// C_XOR/D///      x117y79     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1615_1 ( .OUT(na1615_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na264_1), .IN6(na713_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1615_2 ( .OUT(na1615_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1615_1_i) );
// C_///XOR/D      x113y94     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1616_4 ( .OUT(na1616_2_i), .IN1(1'b0), .IN2(na714_1), .IN3(1'b0), .IN4(na277_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1616_5 ( .OUT(na1616_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1616_2_i) );
// C_XOR/D///      x116y64     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1617_1 ( .OUT(na1617_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na287_1), .IN8(na715_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1617_2 ( .OUT(na1617_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1617_1_i) );
// C_///XOR/D      x93y65     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1618_4 ( .OUT(na1618_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na295_1), .IN4(na716_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1618_5 ( .OUT(na1618_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1618_2_i) );
// C_XOR////D      x82y67     80'hC0_EC18_00_0000_0666_AC03
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1619_1 ( .OUT(na1619_1), .IN1(1'b0), .IN2(~na717_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na303_2), .IN7(na301_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1619_5 ( .OUT(na1619_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1619_1) );
// C_XOR////D      x86y60     80'hC0_EC18_00_0000_0666_60C0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1620_1 ( .OUT(na1620_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na718_1), .IN5(1'b0), .IN6(1'b0), .IN7(na301_2), .IN8(na310_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1620_5 ( .OUT(na1620_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1620_1) );
// C_///XOR/D      x117y61     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1621_4 ( .OUT(na1621_2_i), .IN1(na315_1), .IN2(1'b0), .IN3(1'b0), .IN4(na719_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1621_5 ( .OUT(na1621_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1621_2_i) );
// C_XOR////D      x85y87     80'hC0_EC18_00_0000_0666_0C06
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1622_1 ( .OUT(na1622_1), .IN1(na720_1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na855_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1622_5 ( .OUT(na1622_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1622_1) );
// C_///XOR/D      x105y92     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1623_4 ( .OUT(na1623_2_i), .IN1(na721_1), .IN2(na862_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1623_5 ( .OUT(na1623_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1623_2_i) );
// C_XOR////D      x96y96     80'hC0_EC18_00_0000_0666_065C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1624_1 ( .OUT(na1624_1), .IN1(1'b0), .IN2(na722_1), .IN3(~na874_1), .IN4(1'b0), .IN5(na872_1), .IN6(na873_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1624_5 ( .OUT(na1624_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1624_1) );
// C_XOR/D///      x113y73     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1625_1 ( .OUT(na1625_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na877_1), .IN7(1'b0), .IN8(na723_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1625_2 ( .OUT(na1625_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1625_1_i) );
// C_XOR/D///      x97y78     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1626_1 ( .OUT(na1626_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na724_1), .IN8(na883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1626_2 ( .OUT(na1626_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1626_1_i) );
// C_XOR////D      x81y80     80'hC0_EC18_00_0000_0666_AC06
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1627_1 ( .OUT(na1627_1), .IN1(~na875_1), .IN2(~na725_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na817_1), .IN7(na888_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1627_5 ( .OUT(na1627_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1627_1) );
// C_XOR////D      x84y67     80'hC0_EC18_00_0000_0666_6005
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1628_1 ( .OUT(na1628_1), .IN1(~na726_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na888_1), .IN8(na864_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1628_5 ( .OUT(na1628_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1628_1) );
// C_XOR////D      x87y61     80'hC0_EC18_00_0000_0666_AA0C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1629_1 ( .OUT(na1629_1), .IN1(1'b0), .IN2(na727_1), .IN3(1'b0), .IN4(1'b0), .IN5(na893_2), .IN6(1'b0), .IN7(na888_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1629_5 ( .OUT(na1629_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1629_1) );
// C_XOR/D///      x134y100     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1630_1 ( .OUT(na1630_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na728_1), .IN8(na895_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1630_2 ( .OUT(na1630_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1630_1_i) );
// C_///XOR/D      x132y101     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1631_4 ( .OUT(na1631_2_i), .IN1(1'b0), .IN2(na729_1), .IN3(na4285_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1631_5 ( .OUT(na1631_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1631_2_i) );
// C_XOR////D      x135y101     80'hC0_EC18_00_0000_0666_AC90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1632_1 ( .OUT(na1632_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na952_1), .IN4(na730_1), .IN5(1'b0), .IN6(na950_1), .IN7(na951_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1632_5 ( .OUT(na1632_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1632_1) );
// C_XOR////D      x137y99     80'hC0_EC18_00_0000_0666_6006
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1633_1 ( .OUT(na1633_1), .IN1(~na957_2), .IN2(~na731_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na952_1), .IN8(na956_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1633_5 ( .OUT(na1633_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1633_1) );
// C_///XOR/D      x137y93     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1634_4 ( .OUT(na1634_2_i), .IN1(1'b0), .IN2(na732_1), .IN3(na962_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1634_5 ( .OUT(na1634_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1634_2_i) );
// C_///XOR/D      x131y89     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1635_4 ( .OUT(na1635_2_i), .IN1(1'b0), .IN2(na733_1), .IN3(1'b0), .IN4(na4287_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1635_5 ( .OUT(na1635_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1635_2_i) );
// C_XOR////D      x102y65     80'hC0_EC18_00_0000_0666_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1636_1 ( .OUT(na1636_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na968_1), .IN7(1'b0), .IN8(na734_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1636_5 ( .OUT(na1636_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1636_1) );
// C_XOR/D///      x142y72     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1637_1 ( .OUT(na1637_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na970_1), .IN6(1'b0), .IN7(1'b0), .IN8(na735_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1637_2 ( .OUT(na1637_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1637_1_i) );
// C_XOR////D      x114y100     80'hC0_EC18_00_0000_0666_0630
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1638_1 ( .OUT(na1638_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(~na736_1), .IN5(na1014_1), .IN6(na973_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1638_5 ( .OUT(na1638_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1638_1) );
// C_XOR////D      x115y99     80'hC0_EC18_00_0000_0666_CA0C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1639_1 ( .OUT(na1639_1), .IN1(1'b0), .IN2(na737_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1019_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1022_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1639_5 ( .OUT(na1639_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1639_1) );
// C_XOR////D      x117y102     80'hC0_EC18_00_0000_0666_CC5C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1640_1 ( .OUT(na1640_1), .IN1(1'b0), .IN2(na738_1), .IN3(~na1033_1), .IN4(1'b0), .IN5(1'b0), .IN6(na973_1), .IN7(1'b0), .IN8(na1031_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1640_5 ( .OUT(na1640_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1640_1) );
// C_XOR////D      x113y99     80'hC0_EC18_00_0000_0666_AC3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1641_1 ( .OUT(na1641_1), .IN1(na739_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1036_1), .IN5(1'b0), .IN6(na973_1), .IN7(na1033_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1641_5 ( .OUT(na1641_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1641_1) );
// C_XOR////D      x114y97     80'hC0_EC18_00_0000_0666_630C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1642_1 ( .OUT(na1642_1), .IN1(1'b0), .IN2(na740_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_2), .IN7(na1033_1),
                      .IN8(na1036_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1642_5 ( .OUT(na1642_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1642_1) );
// C_XOR////D      x93y96     80'hC0_EC18_00_0000_0666_AC09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1643_1 ( .OUT(na1643_1), .IN1(~na1026_1), .IN2(na741_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1046_1), .IN7(na1047_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1643_5 ( .OUT(na1643_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1643_1) );
// C_///XOR/D      x108y71     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1644_4 ( .OUT(na1644_2_i), .IN1(na742_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1049_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1644_5 ( .OUT(na1644_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1644_2_i) );
// C_XOR/D///      x113y71     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1645_1 ( .OUT(na1645_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na743_1), .IN7(na1051_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1645_2 ( .OUT(na1645_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1645_1_i) );
// C_XOR/D///      x91y87     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1646_1 ( .OUT(na1646_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na744_1), .IN7(na1614_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1646_2 ( .OUT(na1646_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1646_1_i) );
// C_///XOR/D      x117y79     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1647_4 ( .OUT(na1647_2_i), .IN1(na264_1), .IN2(na713_1), .IN3(na745_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1647_5 ( .OUT(na1647_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1647_2_i) );
// C_XOR/D///      x117y90     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1648_1 ( .OUT(na1648_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na746_1), .IN6(na714_1), .IN7(1'b0), .IN8(na277_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1648_2 ( .OUT(na1648_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1648_1_i) );
// C_///XOR/D      x119y61     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1649_4 ( .OUT(na1649_2_i), .IN1(na747_1), .IN2(1'b0), .IN3(na287_1), .IN4(na715_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1649_5 ( .OUT(na1649_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1649_2_i) );
// C_XOR/D///      x95y66     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1650_1 ( .OUT(na1650_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na748_1), .IN7(na295_1), .IN8(na716_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1650_2 ( .OUT(na1650_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1650_1_i) );
// C_XOR/D///      x81y69     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1651_1 ( .OUT(na1651_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1619_1), .IN8(na749_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1651_2 ( .OUT(na1651_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1651_1_i) );
// C_///XOR/D      x89y61     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1652_4 ( .OUT(na1652_2_i), .IN1(na750_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1620_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1652_5 ( .OUT(na1652_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1652_2_i) );
// C_///XOR/D      x107y61     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1653_4 ( .OUT(na1653_2_i), .IN1(na315_1), .IN2(1'b0), .IN3(na751_1), .IN4(na719_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1653_5 ( .OUT(na1653_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1653_2_i) );
// C_///XOR/D      x81y85     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1654_4 ( .OUT(na1654_2_i), .IN1(na1622_1), .IN2(1'b0), .IN3(na752_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1654_5 ( .OUT(na1654_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1654_2_i) );
// C_XOR/D///      x109y91     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1655_1 ( .OUT(na1655_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na721_1), .IN6(na862_1), .IN7(na753_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1655_2 ( .OUT(na1655_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1655_1_i) );
// C_///XOR/D      x99y96     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1656_4 ( .OUT(na1656_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na754_1), .IN4(na1624_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1656_5 ( .OUT(na1656_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1656_2_i) );
// C_XOR////D      x95y84     80'hC0_EC18_00_0000_0666_CAC5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1657_1 ( .OUT(na1657_1), .IN1(~na755_1), .IN2(1'b0), .IN3(1'b0), .IN4(na723_1), .IN5(na872_1), .IN6(1'b0), .IN7(1'b0), .IN8(na878_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1657_5 ( .OUT(na1657_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1657_1) );
// C_XOR////D      x91y83     80'hC0_EC18_00_0000_0666_CC55
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1658_1 ( .OUT(na1658_1), .IN1(~na756_1), .IN2(1'b0), .IN3(~na724_1), .IN4(1'b0), .IN5(1'b0), .IN6(na884_2), .IN7(1'b0), .IN8(na878_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1658_5 ( .OUT(na1658_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1658_1) );
// C_XOR/D///      x83y78     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1659_1 ( .OUT(na1659_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1627_1), .IN7(na757_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1659_2 ( .OUT(na1659_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1659_1_i) );
// C_XOR/D///      x83y65     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1660_1 ( .OUT(na1660_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na758_1), .IN7(na1628_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1660_2 ( .OUT(na1660_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1660_1_i) );
// C_XOR/D///      x87y63     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1661_1 ( .OUT(na1661_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1629_1), .IN6(1'b0), .IN7(1'b0), .IN8(na759_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1661_2 ( .OUT(na1661_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1661_1_i) );
// C_XOR/D///      x128y99     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1662_1 ( .OUT(na1662_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na760_1), .IN6(1'b0), .IN7(na728_1), .IN8(na895_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1662_2 ( .OUT(na1662_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1662_1_i) );
// C_///XOR/D      x131y102     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1663_4 ( .OUT(na1663_2_i), .IN1(1'b0), .IN2(na729_1), .IN3(na4285_2), .IN4(na761_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1663_5 ( .OUT(na1663_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1663_2_i) );
// C_///XOR/D      x135y97     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1664_4 ( .OUT(na1664_2_i), .IN1(na1632_1), .IN2(na762_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1664_5 ( .OUT(na1664_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1664_2_i) );
// C_XOR/D///      x134y95     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1665_1 ( .OUT(na1665_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1633_1), .IN6(1'b0), .IN7(1'b0), .IN8(na763_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1665_2 ( .OUT(na1665_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1665_1_i) );
// C_XOR////D      x135y92     80'hC0_EC18_00_0000_0666_AA3C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1666_1 ( .OUT(na1666_1), .IN1(1'b0), .IN2(na732_1), .IN3(1'b0), .IN4(~na764_1), .IN5(na963_1), .IN6(1'b0), .IN7(na952_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1666_5 ( .OUT(na1666_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1666_1) );
// C_XOR////D      x124y93     80'hC0_EC18_00_0000_0666_0AA6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1667_1 ( .OUT(na1667_1), .IN1(~na765_1), .IN2(~na733_1), .IN3(na966_2), .IN4(1'b0), .IN5(na963_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1667_5 ( .OUT(na1667_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1667_1) );
// C_XOR/D///      x101y61     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1668_1 ( .OUT(na1668_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na766_1), .IN7(na1636_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1668_2 ( .OUT(na1668_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1668_1_i) );
// C_XOR////D      x131y80     80'hC0_EC18_00_0000_0666_AA35
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1669_1 ( .OUT(na1669_1), .IN1(~na767_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na735_1), .IN5(na963_1), .IN6(1'b0), .IN7(na951_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1669_5 ( .OUT(na1669_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1669_1) );
// C_///XOR/D      x115y102     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1670_4 ( .OUT(na1670_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na768_1), .IN4(na1638_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1670_5 ( .OUT(na1670_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1670_2_i) );
// C_///XOR/D      x113y101     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1671_4 ( .OUT(na1671_2_i), .IN1(na1639_1), .IN2(1'b0), .IN3(na769_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1671_5 ( .OUT(na1671_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1671_2_i) );
// C_///XOR/D      x121y102     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1672_4 ( .OUT(na1672_2_i), .IN1(1'b0), .IN2(na1640_1), .IN3(na770_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1672_5 ( .OUT(na1672_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1672_2_i) );
// C_XOR/D///      x101y93     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1673_1 ( .OUT(na1673_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1641_1), .IN6(1'b0), .IN7(1'b0), .IN8(na771_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1673_2 ( .OUT(na1673_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1673_1_i) );
// C_///XOR/D      x97y94     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1674_4 ( .OUT(na1674_2_i), .IN1(na772_1), .IN2(1'b0), .IN3(na1642_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1674_5 ( .OUT(na1674_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1674_2_i) );
// C_XOR/D///      x91y98     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1675_1 ( .OUT(na1675_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na773_1), .IN6(na1643_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1675_2 ( .OUT(na1675_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1675_1_i) );
// C_XOR////D      x89y77     80'hC0_EC18_00_0000_0666_A0A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1676_1 ( .OUT(na1676_1), .IN1(~na742_1), .IN2(~na774_1), .IN3(na1047_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1023_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1676_5 ( .OUT(na1676_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1676_1) );
// C_XOR////D      x91y77     80'hC0_EC18_00_0000_0666_630C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1677_1 ( .OUT(na1677_1), .IN1(1'b0), .IN2(na743_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na775_1), .IN7(na1047_1), .IN8(na1022_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1677_5 ( .OUT(na1677_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1677_1) );
// C_XOR/D///      x91y90     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1678_1 ( .OUT(na1678_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na744_1), .IN7(na1614_1), .IN8(na776_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1678_2 ( .OUT(na1678_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1678_1_i) );
// C_XOR/D///      x117y81     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1679_1 ( .OUT(na1679_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na264_1), .IN6(~na713_1), .IN7(~na745_1),
                      .IN8(na777_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1679_2 ( .OUT(na1679_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1679_1_i) );
// C_///XOR/D      x116y90     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1680_4 ( .OUT(na1680_2_i), .IN1(~na746_1), .IN2(~na714_1), .IN3(na778_1), .IN4(na277_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1680_5 ( .OUT(na1680_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1680_2_i) );
// C_XOR/D///      x115y61     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1681_1 ( .OUT(na1681_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na747_1), .IN6(na779_1), .IN7(na287_1),
                      .IN8(~na715_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1681_2 ( .OUT(na1681_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1681_1_i) );
// C_///XOR/D      x93y67     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1682_4 ( .OUT(na1682_2_i), .IN1(na4193_2), .IN2(~na748_1), .IN3(na780_1), .IN4(~na716_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1682_5 ( .OUT(na1682_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1682_2_i) );
// C_///XOR/D      x81y72     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1683_4 ( .OUT(na1683_2_i), .IN1(1'b0), .IN2(na781_1), .IN3(na1619_1), .IN4(na749_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1683_5 ( .OUT(na1683_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1683_2_i) );
// C_XOR/D///      x90y60     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1684_1 ( .OUT(na1684_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na750_1), .IN6(na782_1), .IN7(1'b0), .IN8(na1620_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1684_2 ( .OUT(na1684_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1684_1_i) );
// C_///XOR/D      x111y63     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1685_4 ( .OUT(na1685_2_i), .IN1(na315_1), .IN2(na783_1), .IN3(~na751_1), .IN4(~na719_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1685_5 ( .OUT(na1685_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1685_2_i) );
// C_///XOR/D      x91y90     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1686_4 ( .OUT(na1686_2_i), .IN1(na1622_1), .IN2(1'b0), .IN3(na752_1), .IN4(na784_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1686_5 ( .OUT(na1686_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1686_2_i) );
// C_XOR/D///      x107y91     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1687_1 ( .OUT(na1687_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na721_1), .IN6(na862_1), .IN7(~na753_1),
                      .IN8(na785_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1687_2 ( .OUT(na1687_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1687_1_i) );
// C_XOR/D///      x98y93     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1688_1 ( .OUT(na1688_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na786_1), .IN7(na754_1), .IN8(na1624_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1688_2 ( .OUT(na1688_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1688_1_i) );
// C_///XOR/D      x97y79     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1689_4 ( .OUT(na1689_2_i), .IN1(1'b0), .IN2(na1657_1), .IN3(1'b0), .IN4(na787_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1689_5 ( .OUT(na1689_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1689_2_i) );
// C_XOR/D///      x93y84     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1690_1 ( .OUT(na1690_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1658_1), .IN6(1'b0), .IN7(na788_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1690_2 ( .OUT(na1690_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1690_1_i) );
// C_///XOR/D      x84y75     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1691_4 ( .OUT(na1691_2_i), .IN1(1'b0), .IN2(na1627_1), .IN3(na757_1), .IN4(na789_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1691_5 ( .OUT(na1691_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1691_2_i) );
// C_XOR/D///      x85y66     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1692_1 ( .OUT(na1692_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na758_1), .IN7(na1628_1), .IN8(na790_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1692_2 ( .OUT(na1692_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1692_1_i) );
// C_///XOR/D      x91y63     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1693_4 ( .OUT(na1693_2_i), .IN1(na1629_1), .IN2(1'b0), .IN3(na791_1), .IN4(na759_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1693_5 ( .OUT(na1693_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1693_2_i) );
// C_XOR/D///      x130y97     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1694_1 ( .OUT(na1694_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na760_1), .IN6(na792_1), .IN7(~na728_1),
                      .IN8(na895_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1694_2 ( .OUT(na1694_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1694_1_i) );
// C_///XOR/D      x131y99     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1695_4 ( .OUT(na1695_2_i), .IN1(na940_1), .IN2(~na729_1), .IN3(na793_1), .IN4(~na761_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1695_5 ( .OUT(na1695_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1695_2_i) );
// C_XOR/D///      x133y100     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1696_1 ( .OUT(na1696_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1632_1), .IN6(na762_1), .IN7(na794_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1696_2 ( .OUT(na1696_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1696_1_i) );
// C_XOR/D///      x134y96     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1697_1 ( .OUT(na1697_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1633_1), .IN6(1'b0), .IN7(na795_1), .IN8(na763_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1697_2 ( .OUT(na1697_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1697_1_i) );
// C_///XOR/D      x127y90     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1698_4 ( .OUT(na1698_2_i), .IN1(1'b0), .IN2(na1666_1), .IN3(na796_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1698_5 ( .OUT(na1698_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1698_2_i) );
// C_XOR/D///      x117y89     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1699_1 ( .OUT(na1699_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1667_1), .IN8(na797_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1699_2 ( .OUT(na1699_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1699_1_i) );
// C_XOR/D///      x103y66     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1700_1 ( .OUT(na1700_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na766_1), .IN7(na1636_1), .IN8(na798_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1700_2 ( .OUT(na1700_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1700_1_i) );
// C_///XOR/D      x135y68     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1701_4 ( .OUT(na1701_2_i), .IN1(1'b0), .IN2(na1669_1), .IN3(na799_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1701_5 ( .OUT(na1701_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1701_2_i) );
// C_XOR/D///      x115y97     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1702_1 ( .OUT(na1702_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na800_1), .IN7(na768_1), .IN8(na1638_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1702_2 ( .OUT(na1702_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1702_1_i) );
// C_XOR/D///      x118y100     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1703_1 ( .OUT(na1703_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1639_1), .IN6(na801_1), .IN7(na769_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1703_2 ( .OUT(na1703_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1703_1_i) );
// C_XOR/D///      x120y102     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1704_1 ( .OUT(na1704_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1640_1), .IN7(na770_1), .IN8(na802_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1704_2 ( .OUT(na1704_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1704_1_i) );
// C_///XOR/D      x98y93     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1705_4 ( .OUT(na1705_2_i), .IN1(na1641_1), .IN2(1'b0), .IN3(na803_1), .IN4(na771_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1705_5 ( .OUT(na1705_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1705_2_i) );
// C_XOR/D///      x97y92     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1706_1 ( .OUT(na1706_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na772_1), .IN6(na804_1), .IN7(na1642_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1706_2 ( .OUT(na1706_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1706_1_i) );
// C_///XOR/D      x89y89     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1707_4 ( .OUT(na1707_2_i), .IN1(na773_1), .IN2(na1643_1), .IN3(na805_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1707_5 ( .OUT(na1707_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1707_2_i) );
// C_XOR/D///      x89y69     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1708_1 ( .OUT(na1708_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1676_1), .IN6(1'b0), .IN7(1'b0), .IN8(na806_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1708_2 ( .OUT(na1708_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1708_1_i) );
// C_///XOR/D      x87y70     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1709_4 ( .OUT(na1709_2_i), .IN1(na1677_1), .IN2(na807_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1709_5 ( .OUT(na1709_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1709_2_i) );
// C_///XOR/D      x91y82     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1710_4 ( .OUT(na1710_2_i), .IN1(na592_1), .IN2(~na744_1), .IN3(na1614_1), .IN4(~na776_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1710_5 ( .OUT(na1710_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1710_2_i) );
// C_XOR/D///      x115y83     80'hC0_EC00_00_0000_0666_0693
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1711_1 ( .OUT(na1711_1_i), .IN1(1'b0), .IN2(~na713_1), .IN3(~na745_1), .IN4(na777_1), .IN5(na264_1), .IN6(na593_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1711_2 ( .OUT(na1711_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1711_1_i) );
// C_XOR/D///      x115y89     80'hC0_EC00_00_0000_0666_0A66
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1712_1 ( .OUT(na1712_1_i), .IN1(~na746_1), .IN2(~na714_1), .IN3(na778_1), .IN4(na277_1), .IN5(na594_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1712_2 ( .OUT(na1712_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1712_1_i) );
// C_XOR/D///      x110y65     80'hC0_EC00_00_0000_0666_0C99
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1713_1 ( .OUT(na1713_1_i), .IN1(~na747_1), .IN2(na595_1), .IN3(na287_1), .IN4(~na715_1), .IN5(1'b0), .IN6(na779_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1713_2 ( .OUT(na1713_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1713_1_i) );
// C_XOR/D///      x96y71     80'hC0_EC00_00_0000_0666_AC93
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1714_1 ( .OUT(na1714_1_i), .IN1(1'b0), .IN2(~na748_1), .IN3(na780_1), .IN4(~na716_1), .IN5(1'b0), .IN6(na596_1), .IN7(na295_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1714_2 ( .OUT(na1714_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1714_1_i) );
// C_XOR/D///      x85y73     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1715_1 ( .OUT(na1715_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na597_1), .IN6(~na781_1), .IN7(na1619_1),
                      .IN8(~na749_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1715_2 ( .OUT(na1715_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1715_1_i) );
// C_XOR/D///      x91y63     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1716_1 ( .OUT(na1716_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na750_1), .IN6(~na782_1), .IN7(na598_1),
                      .IN8(na1620_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1716_2 ( .OUT(na1716_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1716_1_i) );
// C_XOR/D///      x99y65     80'hC0_EC00_00_0000_0666_563A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1717_1 ( .OUT(na1717_1_i), .IN1(na599_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na719_1), .IN5(na315_1), .IN6(na783_1), .IN7(~na751_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1717_2 ( .OUT(na1717_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1717_1_i) );
// C_///XOR/D      x91y92     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1718_4 ( .OUT(na1718_2_i), .IN1(na1622_1), .IN2(na600_1), .IN3(~na752_1), .IN4(~na784_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1718_5 ( .OUT(na1718_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1718_2_i) );
// C_XOR/D///      x105y94     80'hC0_EC00_00_0000_0666_0C99
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1719_1 ( .OUT(na1719_1_i), .IN1(~na721_1), .IN2(na862_1), .IN3(~na753_1), .IN4(na785_1), .IN5(1'b0), .IN6(na601_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1719_2 ( .OUT(na1719_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1719_1_i) );
// C_XOR/D///      x105y98     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1720_1 ( .OUT(na1720_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na602_1), .IN6(~na786_1), .IN7(~na754_1),
                      .IN8(na1624_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1720_2 ( .OUT(na1720_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1720_1_i) );
// C_XOR/D///      x103y79     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1721_1 ( .OUT(na1721_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1657_1), .IN7(na603_1), .IN8(na787_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1721_2 ( .OUT(na1721_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1721_1_i) );
// C_///XOR/D      x91y75     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1722_4 ( .OUT(na1722_2_i), .IN1(na1658_1), .IN2(na604_1), .IN3(na788_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1722_5 ( .OUT(na1722_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1722_2_i) );
// C_///XOR/D      x85y73     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1723_4 ( .OUT(na1723_2_i), .IN1(na605_1), .IN2(na1627_1), .IN3(~na757_1), .IN4(~na789_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1723_5 ( .OUT(na1723_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1723_2_i) );
// C_///XOR/D      x86y65     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1724_4 ( .OUT(na1724_2_i), .IN1(na606_1), .IN2(~na758_1), .IN3(na1628_1), .IN4(~na790_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1724_5 ( .OUT(na1724_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1724_2_i) );
// C_XOR/D///      x92y64     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1725_1 ( .OUT(na1725_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1629_1), .IN6(na607_1), .IN7(~na791_1),
                      .IN8(~na759_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1725_2 ( .OUT(na1725_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1725_1_i) );
// C_XOR/D///      x127y99     80'hC0_EC00_00_0000_0666_0C99
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1726_1 ( .OUT(na1726_1_i), .IN1(~na760_1), .IN2(na608_1), .IN3(~na728_1), .IN4(na895_1), .IN5(1'b0), .IN6(na792_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1726_2 ( .OUT(na1726_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1726_1_i) );
// C_XOR/D///      x123y104     80'hC0_EC00_00_0000_0666_AC93
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1727_1 ( .OUT(na1727_1_i), .IN1(1'b0), .IN2(~na729_1), .IN3(na793_1), .IN4(~na761_1), .IN5(1'b0), .IN6(na609_1), .IN7(na4285_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1727_2 ( .OUT(na1727_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1727_1_i) );
// C_///XOR/D      x128y97     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1728_4 ( .OUT(na1728_2_i), .IN1(na1632_1), .IN2(~na762_1), .IN3(~na794_1), .IN4(na610_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1728_5 ( .OUT(na1728_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1728_2_i) );
// C_///XOR/D      x124y94     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1729_4 ( .OUT(na1729_2_i), .IN1(na1633_1), .IN2(na611_1), .IN3(~na795_1), .IN4(~na763_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1729_5 ( .OUT(na1729_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1729_2_i) );
// C_XOR/D///      x120y91     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1730_1 ( .OUT(na1730_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4226_2), .IN6(na1666_1), .IN7(na796_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1730_2 ( .OUT(na1730_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1730_1_i) );
// C_XOR/D///      x112y87     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1731_1 ( .OUT(na1731_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na613_1), .IN6(1'b0), .IN7(na1667_1), .IN8(na797_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1731_2 ( .OUT(na1731_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1731_1_i) );
// C_XOR/D///      x97y66     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1732_1 ( .OUT(na1732_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na614_1), .IN6(~na766_1), .IN7(na1636_1),
                      .IN8(~na798_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1732_2 ( .OUT(na1732_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1732_1_i) );
// C_///XOR/D      x117y67     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1733_4 ( .OUT(na1733_2_i), .IN1(1'b0), .IN2(na1669_1), .IN3(na799_1), .IN4(na615_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1733_5 ( .OUT(na1733_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1733_2_i) );
// C_XOR/D///      x103y95     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1734_1 ( .OUT(na1734_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na584_1), .IN6(~na800_1), .IN7(~na768_1),
                      .IN8(na1638_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1734_2 ( .OUT(na1734_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1734_1_i) );
// C_XOR/D///      x107y95     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1735_1 ( .OUT(na1735_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1639_1), .IN6(~na801_1), .IN7(~na769_1),
                      .IN8(na4220_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1735_2 ( .OUT(na1735_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1735_1_i) );
// C_XOR/D///      x117y97     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1736_1 ( .OUT(na1736_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na586_1), .IN6(na1640_1), .IN7(~na770_1),
                      .IN8(~na802_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1736_2 ( .OUT(na1736_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1736_1_i) );
// C_///XOR/D      x99y85     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1737_4 ( .OUT(na1737_2_i), .IN1(na1641_1), .IN2(na587_1), .IN3(~na803_1), .IN4(~na771_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1737_5 ( .OUT(na1737_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1737_2_i) );
// C_XOR/D///      x101y94     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1738_1 ( .OUT(na1738_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na772_1), .IN6(~na804_1), .IN7(na1642_1),
                      .IN8(na588_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1738_2 ( .OUT(na1738_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1738_1_i) );
// C_XOR/D///      x94y95     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1739_1 ( .OUT(na1739_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na589_1), .IN6(na1643_1), .IN7(~na805_1),
                      .IN8(~na4239_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1739_2 ( .OUT(na1739_1), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1739_1_i) );
// C_///XOR/D      x87y69     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1740_4 ( .OUT(na1740_2_i), .IN1(na1676_1), .IN2(na590_1), .IN3(1'b0), .IN4(na806_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1740_5 ( .OUT(na1740_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1740_2_i) );
// C_///XOR/D      x91y74     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1741_4 ( .OUT(na1741_2_i), .IN1(na1677_1), .IN2(na807_1), .IN3(1'b0), .IN4(na591_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1741_5 ( .OUT(na1741_2), .CLK(1'b0), .EN(1'b0), .SR(na3289_1), .CINY2(na4512_3), .PINY2(~na4512_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1741_2_i) );
// C_XOR////      x141y64     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1742_1 ( .OUT(na1742_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na324_1), .IN6(na1743_2), .IN7(na316_1), .IN8(~na397_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y62     80'h00_0060_00_0000_0C06_FFA5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1743_4 ( .OUT(na1743_2), .IN1(~na530_1), .IN2(1'b0), .IN3(na467_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y61     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1744_4 ( .OUT(na1744_2), .IN1(na1745_2), .IN2(na1743_2), .IN3(~na333_1), .IN4(~na1746_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y59     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1745_4 ( .OUT(na1745_2), .IN1(na1819_1), .IN2(1'b0), .IN3(~na316_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y64     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1746_1 ( .OUT(na1746_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na476_1), .IN6(1'b0), .IN7(1'b0), .IN8(na405_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x152y66     80'h00_0018_00_0000_0666_06C6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1747_1 ( .OUT(na1747_1), .IN1(na476_1), .IN2(na1824_1), .IN3(1'b0), .IN4(na485_1), .IN5(na342_1), .IN6(na414_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x141y66     80'h00_0018_00_0000_0666_9A69
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1749_1 ( .OUT(na1749_1), .IN1(~na4194_2), .IN2(na423_1), .IN3(~na279_1), .IN4(~na485_1), .IN5(na530_1), .IN6(1'b0), .IN7(na353_1),
                      .IN8(~na494_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y61     80'h00_0018_00_0000_0666_6695
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1751_1 ( .OUT(na1751_1), .IN1(~na1829_1), .IN2(1'b0), .IN3(~na362_1), .IN4(na4195_2), .IN5(na503_1), .IN6(na432_1), .IN7(na4201_2),
                      .IN8(na494_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x132y62     80'h00_0018_00_0000_0666_CA39
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1753_1 ( .OUT(na1753_1), .IN1(~na503_1), .IN2(na512_1), .IN3(1'b0), .IN4(~na1834_1), .IN5(na441_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na371_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y59     80'h00_0018_00_0000_0666_C39C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1755_1 ( .OUT(na1755_1), .IN1(1'b0), .IN2(na512_1), .IN3(na1838_1), .IN4(~na380_1), .IN5(1'b0), .IN6(~na521_1), .IN7(1'b0),
                      .IN8(na449_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y60     80'h00_0018_00_0000_0666_A909
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1757_1 ( .OUT(na1757_1), .IN1(~na530_1), .IN2(na1862_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na4198_2), .IN6(na521_1), .IN7(na458_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y62     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1759_1 ( .OUT(na1759_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1745_2), .IN6(na389_1), .IN7(na467_1), .IN8(~na397_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x148y62     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1760_4 ( .OUT(na1760_2), .IN1(na1745_2), .IN2(~na1761_2), .IN3(~na4361_2), .IN4(na1746_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x145y60     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1761_4 ( .OUT(na1761_2), .IN1(na324_1), .IN2(~na389_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x147y66     80'h00_0018_00_0000_0666_AC93
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1762_1 ( .OUT(na1762_1), .IN1(1'b0), .IN2(~na1824_1), .IN3(na333_1), .IN4(~na485_1), .IN5(1'b0), .IN6(na414_1), .IN7(na279_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x142y62     80'h00_0018_00_0000_0666_A699
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1764_1 ( .OUT(na1764_1), .IN1(~na342_1), .IN2(na389_1), .IN3(~na279_1), .IN4(na494_1), .IN5(na1829_1), .IN6(na423_1), .IN7(na316_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x138y62     80'h00_0018_00_0000_0666_69A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1766_1 ( .OUT(na1766_1), .IN1(~na503_1), .IN2(na432_1), .IN3(na316_1), .IN4(1'b0), .IN5(~na1829_1), .IN6(na389_1), .IN7(na353_1),
                      .IN8(na1834_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x132y61     80'h00_0018_00_0000_0666_AA93
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1768_1 ( .OUT(na1768_1), .IN1(1'b0), .IN2(~na512_1), .IN3(~na1838_1), .IN4(na1834_1), .IN5(na441_1), .IN6(1'b0), .IN7(na362_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x130y59     80'h00_0018_00_0000_0666_CC6C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1770_1 ( .OUT(na1770_1), .IN1(1'b0), .IN2(na1862_1), .IN3(na1838_1), .IN4(na449_1), .IN5(1'b0), .IN6(na521_1), .IN7(1'b0),
                      .IN8(na371_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y59     80'h00_0018_00_0000_0666_A066
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1772_1 ( .OUT(na1772_1), .IN1(~na530_1), .IN2(~na1862_1), .IN3(na458_1), .IN4(na380_1), .IN5(1'b0), .IN6(1'b0), .IN7(na316_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y61     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1774_1 ( .OUT(na1774_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1819_1), .IN6(na1761_2), .IN7(~na467_1),
                      .IN8(na4199_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x148y63     80'h00_0018_00_0000_0666_AC96
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1775_1 ( .OUT(na1775_1), .IN1(na476_1), .IN2(na1824_1), .IN3(~na333_1), .IN4(na397_1), .IN5(1'b0), .IN6(na1761_2), .IN7(na458_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x153y67     80'h00_0018_00_0000_0666_6A60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1777_1 ( .OUT(na1777_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na333_1), .IN4(~na485_1), .IN5(na342_1), .IN6(1'b0), .IN7(na279_1),
                      .IN8(na405_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x145y63     80'h00_0018_00_0000_0666_A699
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1779_1 ( .OUT(na1779_1), .IN1(~na342_1), .IN2(na389_1), .IN3(~na353_1), .IN4(na494_1), .IN5(na1829_1), .IN6(na414_1), .IN7(na458_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x141y61     80'h00_0018_00_0000_0666_9663
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1781_1 ( .OUT(na1781_1), .IN1(1'b0), .IN2(~na423_1), .IN3(na458_1), .IN4(na1834_1), .IN5(na503_1), .IN6(na389_1), .IN7(~na362_1),
                      .IN8(na4197_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y62     80'h00_0018_00_0000_0666_9C5C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1783_1 ( .OUT(na1783_1), .IN1(1'b0), .IN2(na512_1), .IN3(~na1838_1), .IN4(1'b0), .IN5(1'b0), .IN6(na432_1), .IN7(~na362_1),
                      .IN8(na371_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y59     80'h00_0018_00_0000_0666_363C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1784_1 ( .OUT(na1784_1), .IN1(1'b0), .IN2(na1862_1), .IN3(1'b0), .IN4(~na371_1), .IN5(na441_1), .IN6(na521_1), .IN7(1'b0),
                      .IN8(~na380_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x140y60     80'h00_0018_00_0000_0666_3690
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1785_1 ( .OUT(na1785_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na316_1), .IN4(na449_1), .IN5(na530_1), .IN6(na389_1), .IN7(1'b0),
                      .IN8(~na380_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y62     80'h00_0018_00_0000_0666_9AA5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1787_1 ( .OUT(na1787_1), .IN1(~na324_1), .IN2(1'b0), .IN3(na4200_2), .IN4(1'b0), .IN5(na1819_1), .IN6(1'b0), .IN7(na458_1),
                      .IN8(~na397_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x143y64     80'h00_0018_00_0000_0666_6C9C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1789_1 ( .OUT(na1789_1), .IN1(1'b0), .IN2(na1824_1), .IN3(na333_1), .IN4(~na405_1), .IN5(1'b0), .IN6(na1743_2), .IN7(na458_1),
                      .IN8(na397_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x152y71     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1790_4 ( .OUT(na1790_2), .IN1(~na342_1), .IN2(na414_1), .IN3(~na279_1), .IN4(na1746_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y63     80'h00_0018_00_0000_0666_A699
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1791_1 ( .OUT(na1791_1), .IN1(~na530_1), .IN2(na414_1), .IN3(~na353_1), .IN4(na485_1), .IN5(na1829_1), .IN6(na423_1), .IN7(na458_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x137y64     80'h00_0018_00_0000_0666_6963
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1793_1 ( .OUT(na1793_1), .IN1(1'b0), .IN2(~na423_1), .IN3(na458_1), .IN4(na1834_1), .IN5(na530_1), .IN6(~na432_1), .IN7(na362_1),
                      .IN8(na494_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x131y61     80'h00_0018_00_0000_0666_C655
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1795_1 ( .OUT(na1795_1), .IN1(~na441_1), .IN2(1'b0), .IN3(~na1838_1), .IN4(1'b0), .IN5(na503_1), .IN6(na432_1), .IN7(1'b0),
                      .IN8(na371_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y61     80'h00_0018_00_0000_0666_363C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1797_1 ( .OUT(na1797_1), .IN1(1'b0), .IN2(na512_1), .IN3(1'b0), .IN4(~na449_1), .IN5(na441_1), .IN6(na1862_1), .IN7(1'b0),
                      .IN8(~na380_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x139y60     80'h00_0018_00_0000_0666_A363
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1798_1 ( .OUT(na1798_1), .IN1(1'b0), .IN2(~na521_1), .IN3(na316_1), .IN4(na449_1), .IN5(1'b0), .IN6(~na389_1), .IN7(na458_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y94     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1810_1 ( .OUT(na1810_1), .IN1(1'b1), .IN2(na4432_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1160_1), .IN8(na4106_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x81y93     80'h00_0018_00_0000_0666_3FCB
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1811_1 ( .OUT(na1811_1), .IN1(~na3470_2), .IN2(na227_1), .IN3(1'b1), .IN4(~na1810_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na221_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x91y93     80'h00_0018_00_0040_0A74_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1812_1 ( .OUT(na1812_1), .IN1(1'b1), .IN2(~na4319_2), .IN3(na1160_1), .IN4(1'b1), .IN5(na4316_2), .IN6(na4108_1), .IN7(~na225_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x90y97     80'h00_0018_00_0000_0C66_5700
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1813_1 ( .OUT(na1813_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4109_2), .IN6(na1151_1), .IN7(na233_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x81y94     80'h00_0018_00_0000_0666_5FDA
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1814_1 ( .OUT(na1814_1), .IN1(~na1812_1), .IN2(1'b1), .IN3(na4180_2), .IN4(~na4106_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1813_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y80     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1816_1 ( .OUT(na1816_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na214_2), .IN8(~na2918_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x141y68     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1817_1 ( .OUT(na1817_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na261_2), .IN7(na4114_1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x134y74     80'h00_0018_00_0040_0C43_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1818_1 ( .OUT(na1818_1), .IN1(na4115_1), .IN2(na263_1), .IN3(1'b1), .IN4(1'b0), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x141y65     80'h40_E800_00_0040_0C5A_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1819_1 ( .OUT(na1819_1_i), .IN1(1'b1), .IN2(na4116_2), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(na1817_1), .IN7(1'b1),
                      .IN8(~na1818_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1819_2 ( .OUT(na1819_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1819_1_i) );
// C_MX4b////      x130y78     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1821_1 ( .OUT(na1821_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na4191_2),
                      .IN8(~na2919_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x142y73     80'h00_0060_00_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1822_4 ( .OUT(na1822_2), .IN1(1'b0), .IN2(~na274_1), .IN3(na4119_1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x137y73     80'h00_0018_00_0040_0C43_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1823_1 ( .OUT(na1823_1), .IN1(na4120_1), .IN2(na276_2), .IN3(1'b1), .IN4(1'b0), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x145y66     80'h40_E800_00_0040_0C3C_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1824_1 ( .OUT(na1824_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4121_2), .IN4(na1451_2), .IN5(~na1823_1), .IN6(1'b1), .IN7(na1822_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1824_2 ( .OUT(na1824_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1824_1_i) );
// C_MX4b////      x126y71     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1826_1 ( .OUT(na1826_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na287_2), .IN8(~na2921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x140y65     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1827_1 ( .OUT(na1827_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na292_2), .IN7(na4124_1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x135y69     80'h00_0018_00_0040_0C2C_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1828_1 ( .OUT(na1828_1), .IN1(1'b0), .IN2(1'b1), .IN3(na294_2), .IN4(na4125_1), .IN5(~na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x133y63     80'h40_E800_00_0040_0C3C_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1829_1 ( .OUT(na1829_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4126_1), .IN4(na1451_2), .IN5(~na1828_1), .IN6(1'b1), .IN7(na1827_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1829_2 ( .OUT(na1829_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1829_1_i) );
// C_MX4b////      x122y71     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1831_1 ( .OUT(na1831_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(~na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na295_2), .IN8(~na2922_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x137y66     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1832_1 ( .OUT(na1832_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na297_1), .IN7(na4129_2), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x132y69     80'h00_0018_00_0040_0C43_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1833_1 ( .OUT(na1833_1), .IN1(na4130_1), .IN2(na299_2), .IN3(1'b1), .IN4(1'b0), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x130y62     80'h40_E800_00_0040_0C5A_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1834_1 ( .OUT(na1834_1_i), .IN1(1'b1), .IN2(na4131_1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(na1832_1), .IN7(~na1833_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1834_2 ( .OUT(na1834_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1834_1_i) );
// C_///ORAND/      x123y66     80'h00_0060_00_0000_0C08_FF3D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1835_4 ( .OUT(na1835_2), .IN1(~na307_1), .IN2(na4133_1), .IN3(1'b0), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x121y69     80'h00_0018_00_0040_0C1C_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1836_1 ( .OUT(na1836_1), .IN1(1'b1), .IN2(1'b0), .IN3(na4134_1), .IN4(na308_1), .IN5(na21_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x125y64     80'h00_0018_00_0040_0C71_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1837_1 ( .OUT(na1837_1), .IN1(~na300_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b0), .IN5(~na1836_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x128y61     80'h40_E800_00_0000_0788_FCE3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1838_1 ( .OUT(na1838_1_i), .IN1(1'b0), .IN2(~na1835_2), .IN3(na304_1), .IN4(na1451_2), .IN5(1'b0), .IN6(na1837_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1838_2 ( .OUT(na1838_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1838_1_i) );
// C_MX2b////      x123y60     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1839_1 ( .OUT(na1839_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(na309_1), .IN7(1'b0), .IN8(na1993_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x84y102     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1840_4 ( .OUT(na1840_2), .IN1(1'b0), .IN2(1'b0), .IN3(na4138_1), .IN4(~na826_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x84y101     80'h00_0060_00_0000_0C06_FF3E
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1841_4 ( .OUT(na1841_2), .IN1(~na4244_2), .IN2(~na822_2), .IN3(1'b1), .IN4(na1840_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x79y99     80'h00_0018_00_0000_0C66_AEFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1842_1 ( .OUT(na1842_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4242_2), .IN6(~na827_2), .IN7(~na1841_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y101     80'h00_0018_00_0000_0666_0936
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1844_1 ( .OUT(na1844_1), .IN1(na1178_1), .IN2(na4143_2), .IN3(1'b0), .IN4(~na834_1), .IN5(~na4142_2), .IN6(na4143_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x142y102     80'h00_0018_00_0040_0AFA_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1845_1 ( .OUT(na1845_1), .IN1(1'b1), .IN2(na904_1), .IN3(~na901_1), .IN4(1'b1), .IN5(na4271_2), .IN6(~na900_1), .IN7(na4270_2),
                      .IN8(~na899_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x147y98     80'h00_0060_00_0000_0C06_FF3E
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1846_4 ( .OUT(na1846_2), .IN1(~na3753_2), .IN2(~na4275_2), .IN3(1'b1), .IN4(na1845_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x151y102     80'h00_0060_00_0000_0C06_FFEC
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1847_4 ( .OUT(na1847_2), .IN1(1'b1), .IN2(~na1846_2), .IN3(~na901_2), .IN4(~na903_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x139y99     80'h00_0018_00_0040_0AD3_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1848_1 ( .OUT(na1848_1), .IN1(1'b1), .IN2(na4404_2), .IN3(1'b1), .IN4(na4399_2), .IN5(~na3753_1), .IN6(1'b1), .IN7(na1184_1),
                      .IN8(na4272_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x93y97     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1850_1 ( .OUT(na1850_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na982_1), .IN6(na4148_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x94y101     80'h00_0060_00_0000_0C06_FFE5
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1851_4 ( .OUT(na1851_2), .IN1(na1850_1), .IN2(1'b1), .IN3(~na4297_2), .IN4(~na3793_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x95y101     80'h00_0018_00_0000_0C66_AEFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1852_1 ( .OUT(na1852_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na977_2), .IN6(~na4295_2), .IN7(~na1851_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y97     80'h00_0018_00_0040_0A7C_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1853_1 ( .OUT(na1853_1), .IN1(1'b1), .IN2(na979_2), .IN3(1'b1), .IN4(~na3793_2), .IN5(na1200_1), .IN6(na979_1), .IN7(~na4415_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x156y79     80'h00_0018_00_0040_0A90_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1855_1 ( .OUT(na1855_1), .IN1(na10_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4168_2), .IN5(na961_1), .IN6(1'b0), .IN7(1'b0), .IN8(na1120_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x151y75     80'h00_0018_00_0000_0888_2222
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1856_1 ( .OUT(na1856_1), .IN1(na1283_1), .IN2(~na1277_1), .IN3(na1280_1), .IN4(~na4006_1), .IN5(na4003_2), .IN6(~na1277_2),
                      .IN7(na4005_2), .IN8(~na4006_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x148y68     80'h40_E800_00_0000_0388_7AFF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1857_1 ( .OUT(na1857_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1856_1), .IN6(1'b0), .IN7(~na1855_1), .IN8(~na1223_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1857_2 ( .OUT(na1857_1), .CLK(1'b0), .EN(na7_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1857_1_i) );
// C_MX2b////      x122y66     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1858_1 ( .OUT(na1858_1), .IN1(1'b1), .IN2(~na1859_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1387_2), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/DST///      x121y70     80'h60_BC00_00_0040_0AE1_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1859_1 ( .OUT(na1859_1_i), .IN1(~na1331_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1332_1), .IN5(1'b1), .IN6(na4433_2), .IN7(na4155_1),
                      .IN8(na4154_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0000)) 
           _a1859_2 ( .OUT(na1859_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1859_1_i) );
// C_MX2b////      x125y62     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1861_1 ( .OUT(na1861_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b0), .IN6(na4157_2), .IN7(1'b0), .IN8(na314_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x127y60     80'h40_E800_00_0000_0788_FC5B
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1862_1 ( .OUT(na1862_1_i), .IN1(na21_2), .IN2(~na1839_1), .IN3(~na312_1), .IN4(1'b0), .IN5(1'b0), .IN6(na1861_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1862_2 ( .OUT(na1862_1), .CLK(1'b0), .EN(na552_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1862_1_i) );
// C_ADDF2///ADDF2/      x143y84     80'h00_0078_00_0020_0C66_3503
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1864_1 ( .OUT(na1864_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1253_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1219_1),
                      .CINX(1'b0), .CINY1(na1871_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1864_4 ( .OUT(na1864_2), .COUTY1(na1864_4), .IN1(1'b1), .IN2(~na1265_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1253_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(~na1219_1), .CINX(1'b0), .CINY1(na1871_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y85     80'h00_0078_00_0020_0C66_3003
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1866_1 ( .OUT(na1866_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na1857_1),
                      .CINX(1'b0), .CINY1(na1864_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1866_4 ( .OUT(na1866_2), .COUTY1(na1866_4), .IN1(1'b1), .IN2(~na1286_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b1), .IN8(~na1857_1), .CINX(1'b0), .CINY1(na1864_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y86     80'h00_0078_00_0020_0C66_5050
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1868_1 ( .OUT(na1868_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1297_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1866_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1868_4 ( .OUT(na1868_2), .COUTY1(na1868_4), .IN1(1'b0), .IN2(1'b0), .IN3(~na1308_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(~na1297_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na1866_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x143y87     80'h00_0018_00_0010_0666_0005
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1870_1 ( .OUT(na1870_1), .COUTY1(na1870_4), .IN1(~na1319_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1868_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x143y83     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1871_2 ( .OUT(na1871_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1871_6 ( .COUTY1(na1871_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1871_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x90y91     80'h00_0078_00_0020_0C66_AA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1872_1 ( .OUT(na1872_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3_2), .IN6(1'b1), .IN7(na2_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1877_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1872_4 ( .OUT(na1872_2), .COUTY1(na1872_4), .IN1(na3_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3_2), .IN6(1'b1), .IN7(na2_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1877_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y92     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1874_1 ( .OUT(na1874_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na5_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1872_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1874_4 ( .OUT(na1874_2), .COUTY1(na1874_4), .IN1(1'b1), .IN2(na5_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na5_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na1872_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x90y93     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1876_1 ( .OUT(na1876_1), .IN1(na6_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1874_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x90y90     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1877_2 ( .OUT(na1877_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1877_6 ( .COUTY1(na1877_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1877_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x145y83     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1878_1 ( .OUT(na1878_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na10_2), .IN6(1'b1), .IN7(1'b1), .IN8(na9_2),
                      .CINX(1'b0), .CINY1(na1882_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1878_4 ( .OUT(na1878_2), .COUTY1(na1878_4), .IN1(na10_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na10_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na9_2), .CINX(1'b0), .CINY1(na1882_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x145y84     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1880_1 ( .OUT(na1880_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na12_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1878_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1880_4 ( .OUT(na1880_2), .IN1(1'b1), .IN2(na12_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na12_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1878_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x145y82     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1882_2 ( .OUT(na1882_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1882_6 ( .COUTY1(na1882_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1882_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x128y75     80'h00_0078_00_0020_0C66_AC0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1883_1 ( .OUT(na1883_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1333_2), .IN7(na4342_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1886_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1883_4 ( .OUT(na1883_2), .COUTY1(na1883_4), .IN1(na1335_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1333_2),
                      .IN7(na4342_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1886_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x128y76     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1885_1 ( .OUT(na1885_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1336_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1883_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x128y74     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1886_2 ( .OUT(na1886_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1886_6 ( .COUTY1(na1886_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1886_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x89y71     80'h00_0078_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1888_1 ( .OUT(na1888_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1351_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1346_1),
                      .CINX(1'b0), .CINY1(na1897_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1888_4 ( .OUT(na1888_2), .COUTY1(na1888_4), .IN1(1'b1), .IN2(na1355_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1351_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na1346_1), .CINX(1'b0), .CINY1(na1897_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y72     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1890_1 ( .OUT(na1890_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1353_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1888_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1890_4 ( .OUT(na1890_2), .COUTY1(na1890_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1359_2), .IN4(1'b1), .IN5(1'b1), .IN6(na1353_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1888_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y73     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1892_1 ( .OUT(na1892_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1355_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1890_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1892_4 ( .OUT(na1892_2), .COUTY1(na1892_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1356_2), .IN5(1'b1), .IN6(na1355_1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1890_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y74     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1894_1 ( .OUT(na1894_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1357_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1892_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1894_4 ( .OUT(na1894_2), .COUTY1(na1894_4), .IN1(na1358_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1357_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1892_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x89y75     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1896_1 ( .OUT(na1896_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1359_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1894_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1896_4 ( .OUT(na1896_2), .IN1(na1358_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1359_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1894_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x89y70     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1897_2 ( .OUT(na1897_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1897_6 ( .COUTY1(na1897_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1897_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x89y79     80'h00_0078_00_0020_0C66_ACC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1898_1 ( .OUT(na1898_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na4344_2), .IN7(na1343_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1900_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1898_4 ( .OUT(na1898_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1345_1), .IN5(1'b1), .IN6(na4344_2), .IN7(na1343_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1900_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x89y78     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1900_2 ( .OUT(na1900_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1900_6 ( .COUTY1(na1900_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1900_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x143y69     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1902_1 ( .OUT(na1902_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1370_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1376_1),
                      .CINX(1'b0), .CINY1(na1911_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1902_4 ( .OUT(na1902_2), .COUTY1(na1902_4), .IN1(na1377_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1370_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na1376_1), .CINX(1'b0), .CINY1(na1911_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y70     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1904_1 ( .OUT(na1904_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1378_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1902_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1904_4 ( .OUT(na1904_2), .COUTY1(na1904_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1379_1), .IN4(1'b1), .IN5(1'b1), .IN6(na1378_1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1902_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y71     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1906_1 ( .OUT(na1906_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1380_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1904_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1906_4 ( .OUT(na1906_2), .COUTY1(na1906_4), .IN1(na1377_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1380_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1904_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y72     80'h00_0078_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1908_1 ( .OUT(na1908_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1382_2),
                      .CINX(1'b0), .CINY1(na1906_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1908_4 ( .OUT(na1908_2), .COUTY1(na1908_4), .IN1(1'b1), .IN2(na1383_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na1382_2), .CINX(1'b0), .CINY1(na1906_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x143y73     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1910_1 ( .OUT(na1910_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1383_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1908_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1910_4 ( .OUT(na1910_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1379_2), .IN4(1'b1), .IN5(1'b1), .IN6(na1383_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1908_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x143y68     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1911_2 ( .OUT(na1911_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1911_6 ( .COUTY1(na1911_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1911_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x145y76     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1912_1 ( .OUT(na1912_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1216_2), .IN7(na1217_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3296_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1912_4 ( .OUT(na1912_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1217_1), .IN4(1'b1), .IN5(1'b1), .IN6(na1216_2), .IN7(na1217_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3296_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x109y92     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1915_1 ( .OUT(na1915_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3173_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1915_2 ( .OUT(na1915_1), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1915_1_i) );
// C_///AND/D      x125y103     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1916_4 ( .OUT(na1916_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1916_5 ( .OUT(na1916_2), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1916_2_i) );
// C_AND/D///      x122y100     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1917_1 ( .OUT(na1917_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3175_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1917_2 ( .OUT(na1917_1), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1917_1_i) );
// C_///AND/D      x120y79     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1918_4 ( .OUT(na1918_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3176_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1918_5 ( .OUT(na1918_2), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1918_2_i) );
// C_AND/D///      x108y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1919_1 ( .OUT(na1919_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3177_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1919_2 ( .OUT(na1919_1), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1919_1_i) );
// C_///AND/D      x86y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1920_4 ( .OUT(na1920_2_i), .IN1(1'b1), .IN2(na3178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1920_5 ( .OUT(na1920_2), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1920_2_i) );
// C_///AND/D      x103y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1921_4 ( .OUT(na1921_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1921_5 ( .OUT(na1921_2), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1921_2_i) );
// C_AND/D///      x105y62     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1922_1 ( .OUT(na1922_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1922_2 ( .OUT(na1922_1), .CLK(1'b0), .EN(na1388_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1922_1_i) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0000_0010)) 
           _a1923 ( .GLB0(na1923_1), .GLB1(_d3), .GLB2(_d4), .GLB3(_d5), .CLK_FB0(_d6), .CLK_FB1(_d7), .CLK_FB2(_d8), .CLK_FB3(_d9),
                    .CLK0_0(1'b0), .CLK0_90(1'b0), .CLK0_180(1'b0), .CLK0_270(1'b0), .CLK0_BYP(na1_1), .CLK1_0(1'b0), .CLK1_90(1'b0),
                    .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                    .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(1'b0),
                    .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_///AND/D      x99y95     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1924_4 ( .OUT(na1924_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1924_5 ( .OUT(na1924_2), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1924_2_i) );
// C_AND/D///      x123y95     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1925_1 ( .OUT(na1925_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1925_2 ( .OUT(na1925_1), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1925_1_i) );
// C_///AND/D      x119y95     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1926_4 ( .OUT(na1926_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1926_5 ( .OUT(na1926_2), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1926_2_i) );
// C_AND/D///      x113y80     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1927_1 ( .OUT(na1927_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1927_2 ( .OUT(na1927_1), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1927_1_i) );
// C_///AND/D      x101y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1928_4 ( .OUT(na1928_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1928_5 ( .OUT(na1928_2), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1928_2_i) );
// C_AND/D///      x83y74     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1929_1 ( .OUT(na1929_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1929_2 ( .OUT(na1929_1), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1929_1_i) );
// C_///AND/D      x104y66     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1930_4 ( .OUT(na1930_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1930_5 ( .OUT(na1930_2), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1930_2_i) );
// C_AND/D///      x96y63     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1931_1 ( .OUT(na1931_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1931_2 ( .OUT(na1931_1), .CLK(1'b0), .EN(na1480_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1931_1_i) );
// C_///AND/D      x124y90     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1961_4 ( .OUT(na1961_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1961_5 ( .OUT(na1961_2), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1961_2_i) );
// C_AND/D///      x127y96     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1962_1 ( .OUT(na1962_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1962_2 ( .OUT(na1962_1), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1962_1_i) );
// C_///AND/D      x131y95     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1963_4 ( .OUT(na1963_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1963_5 ( .OUT(na1963_2), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1963_2_i) );
// C_AND/D///      x132y83     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1964_1 ( .OUT(na1964_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1964_2 ( .OUT(na1964_1), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1964_1_i) );
// C_///AND/D      x112y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1965_4 ( .OUT(na1965_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1965_5 ( .OUT(na1965_2), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1965_2_i) );
// C_AND/D///      x105y78     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1966_1 ( .OUT(na1966_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1966_2 ( .OUT(na1966_1), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1966_1_i) );
// C_///AND/D      x111y65     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1967_4 ( .OUT(na1967_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1967_5 ( .OUT(na1967_2), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1967_2_i) );
// C_AND/D///      x110y60     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1968_1 ( .OUT(na1968_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1968_2 ( .OUT(na1968_1), .CLK(1'b0), .EN(na1422_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1968_1_i) );
// C_///AND/D      x107y84     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1971_4 ( .OUT(na1971_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1971_5 ( .OUT(na1971_2), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1971_2_i) );
// C_AND/D///      x127y94     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1972_1 ( .OUT(na1972_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1972_2 ( .OUT(na1972_1), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1972_1_i) );
// C_///AND/D      x127y94     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1973_4 ( .OUT(na1973_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1973_5 ( .OUT(na1973_2), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1973_2_i) );
// C_AND/D///      x117y76     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1974_1 ( .OUT(na1974_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1974_2 ( .OUT(na1974_1), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1974_1_i) );
// C_///AND/D      x113y72     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1975_4 ( .OUT(na1975_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1975_5 ( .OUT(na1975_2), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1975_2_i) );
// C_AND/D///      x95y72     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1976_1 ( .OUT(na1976_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1976_2 ( .OUT(na1976_1), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1976_1_i) );
// C_///AND/D      x113y62     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1977_4 ( .OUT(na1977_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1977_5 ( .OUT(na1977_2), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1977_2_i) );
// C_AND/D///      x111y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1978_1 ( .OUT(na1978_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1978_2 ( .OUT(na1978_1), .CLK(1'b0), .EN(na1403_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1978_1_i) );
// C_///AND/D      x103y84     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1979_4 ( .OUT(na1979_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1979_5 ( .OUT(na1979_2), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1979_2_i) );
// C_AND/D///      x123y94     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1980_1 ( .OUT(na1980_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1980_2 ( .OUT(na1980_1), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1980_1_i) );
// C_///AND/D      x123y94     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1981_4 ( .OUT(na1981_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1981_5 ( .OUT(na1981_2), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1981_2_i) );
// C_AND/D///      x115y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1982_1 ( .OUT(na1982_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1982_2 ( .OUT(na1982_1), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1982_1_i) );
// C_///AND/D      x107y74     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1983_4 ( .OUT(na1983_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1983_5 ( .OUT(na1983_2), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1983_2_i) );
// C_///AND/D      x85y68     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1984_4 ( .OUT(na1984_2_i), .IN1(1'b1), .IN2(na3178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1984_5 ( .OUT(na1984_2), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1984_2_i) );
// C_///AND/D      x113y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1985_4 ( .OUT(na1985_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1985_5 ( .OUT(na1985_2), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1985_2_i) );
// C_AND/D///      x109y58     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1986_1 ( .OUT(na1986_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1986_2 ( .OUT(na1986_1), .CLK(1'b0), .EN(na1404_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1986_1_i) );
// C_///AND/D      x107y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1987_4 ( .OUT(na1987_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1987_5 ( .OUT(na1987_2), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1987_2_i) );
// C_AND/D///      x129y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1988_1 ( .OUT(na1988_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1988_2 ( .OUT(na1988_1), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1988_1_i) );
// C_///AND/D      x127y88     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1989_4 ( .OUT(na1989_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1989_5 ( .OUT(na1989_2), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1989_2_i) );
// C_AND/D///      x117y71     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1990_1 ( .OUT(na1990_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1990_2 ( .OUT(na1990_1), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1990_1_i) );
// C_///AND/D      x109y73     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1991_4 ( .OUT(na1991_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1991_5 ( .OUT(na1991_2), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1991_2_i) );
// C_AND/D///      x91y71     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1992_1 ( .OUT(na1992_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1992_2 ( .OUT(na1992_1), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1992_1_i) );
// C_///AND/D      x122y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1993_4 ( .OUT(na1993_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1993_5 ( .OUT(na1993_2), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1993_2_i) );
// C_AND/D///      x120y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1994_1 ( .OUT(na1994_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1994_2 ( .OUT(na1994_1), .CLK(1'b0), .EN(na1406_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1994_1_i) );
// C_///AND/D      x108y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1995_4 ( .OUT(na1995_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1995_5 ( .OUT(na1995_2), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1995_2_i) );
// C_AND/D///      x126y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1996_1 ( .OUT(na1996_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1996_2 ( .OUT(na1996_1), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1996_1_i) );
// C_///AND/D      x122y91     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1997_4 ( .OUT(na1997_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1997_5 ( .OUT(na1997_2), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1997_2_i) );
// C_AND/D///      x112y77     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1998_1 ( .OUT(na1998_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1998_2 ( .OUT(na1998_1), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1998_1_i) );
// C_///AND/D      x110y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1999_4 ( .OUT(na1999_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1999_5 ( .OUT(na1999_2), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1999_2_i) );
// C_AND/D///      x92y77     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2000_1 ( .OUT(na2000_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2000_2 ( .OUT(na2000_1), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2000_1_i) );
// C_///AND/D      x112y61     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2001_4 ( .OUT(na2001_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2001_5 ( .OUT(na2001_2), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2001_2_i) );
// C_AND/D///      x112y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2002_1 ( .OUT(na2002_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2002_2 ( .OUT(na2002_1), .CLK(1'b0), .EN(na1407_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2002_1_i) );
// C_///AND/D      x110y83     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2003_4 ( .OUT(na2003_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2003_5 ( .OUT(na2003_2), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2003_2_i) );
// C_AND/D///      x128y93     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2004_1 ( .OUT(na2004_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2004_2 ( .OUT(na2004_1), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2004_1_i) );
// C_///AND/D      x124y95     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2005_4 ( .OUT(na2005_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2005_5 ( .OUT(na2005_2), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2005_2_i) );
// C_AND/D///      x120y75     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2006_1 ( .OUT(na2006_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2006_2 ( .OUT(na2006_1), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2006_1_i) );
// C_///AND/D      x108y77     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2007_4 ( .OUT(na2007_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2007_5 ( .OUT(na2007_2), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2007_2_i) );
// C_AND/D///      x94y69     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2008_1 ( .OUT(na2008_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2008_2 ( .OUT(na2008_1), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2008_1_i) );
// C_///AND/D      x116y59     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2009_4 ( .OUT(na2009_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2009_5 ( .OUT(na2009_2), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2009_2_i) );
// C_AND/D///      x106y61     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2010_1 ( .OUT(na2010_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2010_2 ( .OUT(na2010_1), .CLK(1'b0), .EN(na1409_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2010_1_i) );
// C_///AND/D      x106y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2011_4 ( .OUT(na2011_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2011_5 ( .OUT(na2011_2), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2011_2_i) );
// C_AND/D///      x122y93     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2012_1 ( .OUT(na2012_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2012_2 ( .OUT(na2012_1), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2012_1_i) );
// C_///AND/D      x122y93     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2013_4 ( .OUT(na2013_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2013_5 ( .OUT(na2013_2), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2013_2_i) );
// C_AND/D///      x114y73     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2014_1 ( .OUT(na2014_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2014_2 ( .OUT(na2014_1), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2014_1_i) );
// C_///AND/D      x106y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2015_4 ( .OUT(na2015_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2015_5 ( .OUT(na2015_2), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2015_2_i) );
// C_AND/D///      x92y73     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2016_1 ( .OUT(na2016_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2016_2 ( .OUT(na2016_1), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2016_1_i) );
// C_///AND/D      x116y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2017_4 ( .OUT(na2017_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2017_5 ( .OUT(na2017_2), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2017_2_i) );
// C_AND/D///      x108y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2018_1 ( .OUT(na2018_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2018_2 ( .OUT(na2018_1), .CLK(1'b0), .EN(na1410_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2018_1_i) );
// C_///AND/D      x114y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2019_4 ( .OUT(na2019_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2019_5 ( .OUT(na2019_2), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2019_2_i) );
// C_AND/D///      x130y89     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2020_1 ( .OUT(na2020_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2020_2 ( .OUT(na2020_1), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2020_1_i) );
// C_///AND/D      x126y87     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2021_4 ( .OUT(na2021_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2021_5 ( .OUT(na2021_2), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2021_2_i) );
// C_AND/D///      x120y71     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2022_1 ( .OUT(na2022_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2022_2 ( .OUT(na2022_1), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2022_1_i) );
// C_///AND/D      x118y71     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2023_4 ( .OUT(na2023_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2023_5 ( .OUT(na2023_2), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2023_2_i) );
// C_AND/D///      x98y73     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2024_1 ( .OUT(na2024_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2024_2 ( .OUT(na2024_1), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2024_1_i) );
// C_///AND/D      x114y59     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2025_4 ( .OUT(na2025_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2025_5 ( .OUT(na2025_2), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2025_2_i) );
// C_AND/D///      x106y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2026_1 ( .OUT(na2026_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2026_2 ( .OUT(na2026_1), .CLK(1'b0), .EN(na1411_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2026_1_i) );
// C_///AND/D      x107y90     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2027_4 ( .OUT(na2027_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2027_5 ( .OUT(na2027_2), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2027_2_i) );
// C_AND/D///      x124y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2028_1 ( .OUT(na2028_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2028_2 ( .OUT(na2028_1), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2028_1_i) );
// C_///AND/D      x125y92     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2029_4 ( .OUT(na2029_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2029_5 ( .OUT(na2029_2), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2029_2_i) );
// C_AND/D///      x115y76     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2030_1 ( .OUT(na2030_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2030_2 ( .OUT(na2030_1), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2030_1_i) );
// C_///AND/D      x107y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2031_4 ( .OUT(na2031_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2031_5 ( .OUT(na2031_2), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2031_2_i) );
// C_AND/D///      x98y75     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2032_1 ( .OUT(na2032_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2032_2 ( .OUT(na2032_1), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2032_1_i) );
// C_///AND/D      x113y64     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2033_4 ( .OUT(na2033_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2033_5 ( .OUT(na2033_2), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2033_2_i) );
// C_AND/D///      x111y60     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2034_1 ( .OUT(na2034_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2034_2 ( .OUT(na2034_1), .CLK(1'b0), .EN(na1412_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2034_1_i) );
// C_///AND/D      x108y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2035_4 ( .OUT(na2035_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2035_5 ( .OUT(na2035_2), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2035_2_i) );
// C_AND/D///      x123y98     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2036_1 ( .OUT(na2036_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2036_2 ( .OUT(na2036_1), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2036_1_i) );
// C_///AND/D      x123y98     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2037_4 ( .OUT(na2037_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2037_5 ( .OUT(na2037_2), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2037_2_i) );
// C_AND/D///      x117y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2038_1 ( .OUT(na2038_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2038_2 ( .OUT(na2038_1), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2038_1_i) );
// C_///AND/D      x108y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2039_4 ( .OUT(na2039_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2039_5 ( .OUT(na2039_2), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2039_2_i) );
// C_AND/D///      x92y71     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2040_1 ( .OUT(na2040_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2040_2 ( .OUT(na2040_1), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2040_1_i) );
// C_///AND/D      x117y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2041_4 ( .OUT(na2041_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2041_5 ( .OUT(na2041_2), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2041_2_i) );
// C_AND/D///      x112y65     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2042_1 ( .OUT(na2042_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2042_2 ( .OUT(na2042_1), .CLK(1'b0), .EN(na1414_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2042_1_i) );
// C_///AND/D      x107y86     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2043_4 ( .OUT(na2043_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2043_5 ( .OUT(na2043_2), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2043_2_i) );
// C_AND/D///      x119y92     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2044_1 ( .OUT(na2044_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2044_2 ( .OUT(na2044_1), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2044_1_i) );
// C_AND/D///      x131y94     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2045_1 ( .OUT(na2045_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3175_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2045_2 ( .OUT(na2045_1), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2045_1_i) );
// C_AND/D///      x113y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2046_1 ( .OUT(na2046_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2046_2 ( .OUT(na2046_1), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2046_1_i) );
// C_///AND/D      x105y72     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2047_4 ( .OUT(na2047_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2047_5 ( .OUT(na2047_2), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2047_2_i) );
// C_AND/D///      x92y75     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2048_1 ( .OUT(na2048_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2048_2 ( .OUT(na2048_1), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2048_1_i) );
// C_///AND/D      x113y58     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2049_4 ( .OUT(na2049_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2049_5 ( .OUT(na2049_2), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2049_2_i) );
// C_AND/D///      x110y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2050_1 ( .OUT(na2050_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2050_2 ( .OUT(na2050_1), .CLK(1'b0), .EN(na1415_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2050_1_i) );
// C_///AND/D      x113y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2051_4 ( .OUT(na2051_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2051_5 ( .OUT(na2051_2), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2051_2_i) );
// C_AND/D///      x125y90     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2052_1 ( .OUT(na2052_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2052_2 ( .OUT(na2052_1), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2052_1_i) );
// C_///AND/D      x123y92     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2053_4 ( .OUT(na2053_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2053_5 ( .OUT(na2053_2), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2053_2_i) );
// C_AND/D///      x117y72     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2054_1 ( .OUT(na2054_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2054_2 ( .OUT(na2054_1), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2054_1_i) );
// C_///AND/D      x117y72     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2055_4 ( .OUT(na2055_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2055_5 ( .OUT(na2055_2), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2055_2_i) );
// C_AND/D///      x99y74     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2056_1 ( .OUT(na2056_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2056_2 ( .OUT(na2056_1), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2056_1_i) );
// C_///AND/D      x111y58     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2057_4 ( .OUT(na2057_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2057_5 ( .OUT(na2057_2), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2057_2_i) );
// C_AND/D///      x107y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2058_1 ( .OUT(na2058_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2058_2 ( .OUT(na2058_1), .CLK(1'b0), .EN(na1416_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2058_1_i) );
// C_///AND/D      x108y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2059_4 ( .OUT(na2059_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2059_5 ( .OUT(na2059_2), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2059_2_i) );
// C_AND/D///      x121y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2060_1 ( .OUT(na2060_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2060_2 ( .OUT(na2060_1), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2060_1_i) );
// C_///AND/D      x122y87     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2061_4 ( .OUT(na2061_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2061_5 ( .OUT(na2061_2), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2061_2_i) );
// C_AND/D///      x118y75     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2062_1 ( .OUT(na2062_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2062_2 ( .OUT(na2062_1), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2062_1_i) );
// C_///AND/D      x112y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2063_4 ( .OUT(na2063_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2063_5 ( .OUT(na2063_2), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2063_2_i) );
// C_AND/D///      x93y79     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2064_1 ( .OUT(na2064_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2064_2 ( .OUT(na2064_1), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2064_1_i) );
// C_///AND/D      x110y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2065_4 ( .OUT(na2065_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2065_5 ( .OUT(na2065_2), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2065_2_i) );
// C_AND/D///      x112y57     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2066_1 ( .OUT(na2066_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2066_2 ( .OUT(na2066_1), .CLK(1'b0), .EN(na1417_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2066_1_i) );
// C_///AND/D      x111y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2067_4 ( .OUT(na2067_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2067_5 ( .OUT(na2067_2), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2067_2_i) );
// C_AND/D///      x132y97     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2068_1 ( .OUT(na2068_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2068_2 ( .OUT(na2068_1), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2068_1_i) );
// C_///AND/D      x126y93     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2069_4 ( .OUT(na2069_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2069_5 ( .OUT(na2069_2), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2069_2_i) );
// C_AND/D///      x118y73     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2070_1 ( .OUT(na2070_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2070_2 ( .OUT(na2070_1), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2070_1_i) );
// C_///AND/D      x111y77     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2071_4 ( .OUT(na2071_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2071_5 ( .OUT(na2071_2), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2071_2_i) );
// C_AND/D///      x91y73     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2072_1 ( .OUT(na2072_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2072_2 ( .OUT(na2072_1), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2072_1_i) );
// C_///AND/D      x118y59     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2073_4 ( .OUT(na2073_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2073_5 ( .OUT(na2073_2), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2073_2_i) );
// C_AND/D///      x109y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2074_1 ( .OUT(na2074_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2074_2 ( .OUT(na2074_1), .CLK(1'b0), .EN(na1425_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2074_1_i) );
// C_///AND/D      x101y95     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2075_4 ( .OUT(na2075_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2075_5 ( .OUT(na2075_2), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2075_2_i) );
// C_AND/D///      x119y99     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2076_1 ( .OUT(na2076_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2076_2 ( .OUT(na2076_1), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2076_1_i) );
// C_///AND/D      x119y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2077_4 ( .OUT(na2077_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2077_5 ( .OUT(na2077_2), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2077_2_i) );
// C_AND/D///      x107y83     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2078_1 ( .OUT(na2078_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2078_2 ( .OUT(na2078_1), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2078_1_i) );
// C_///AND/D      x97y86     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2079_4 ( .OUT(na2079_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2079_5 ( .OUT(na2079_2), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2079_2_i) );
// C_AND/D///      x86y82     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2080_1 ( .OUT(na2080_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2080_2 ( .OUT(na2080_1), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2080_1_i) );
// C_///AND/D      x94y65     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2081_4 ( .OUT(na2081_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2081_5 ( .OUT(na2081_2), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2081_2_i) );
// C_AND/D///      x95y61     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2082_1 ( .OUT(na2082_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2082_2 ( .OUT(na2082_1), .CLK(1'b0), .EN(na1418_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2082_1_i) );
// C_///AND/D      x90y80     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2083_4 ( .OUT(na2083_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2083_5 ( .OUT(na2083_2), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2083_2_i) );
// C_AND/D///      x124y88     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2084_1 ( .OUT(na2084_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2084_2 ( .OUT(na2084_1), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2084_1_i) );
// C_///AND/D      x118y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2085_4 ( .OUT(na2085_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2085_5 ( .OUT(na2085_2), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2085_2_i) );
// C_AND/D///      x110y67     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2086_1 ( .OUT(na2086_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2086_2 ( .OUT(na2086_1), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2086_1_i) );
// C_///AND/D      x95y71     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2087_4 ( .OUT(na2087_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2087_5 ( .OUT(na2087_2), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2087_2_i) );
// C_AND/D///      x86y67     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2088_1 ( .OUT(na2088_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2088_2 ( .OUT(na2088_1), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2088_1_i) );
// C_///AND/D      x107y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2089_4 ( .OUT(na2089_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2089_5 ( .OUT(na2089_2), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2089_2_i) );
// C_AND/D///      x105y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2090_1 ( .OUT(na2090_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2090_2 ( .OUT(na2090_1), .CLK(1'b0), .EN(na1420_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2090_1_i) );
// C_///AND/D      x93y83     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2091_4 ( .OUT(na2091_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2091_5 ( .OUT(na2091_2), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2091_2_i) );
// C_AND/D///      x110y89     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2092_1 ( .OUT(na2092_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2092_2 ( .OUT(na2092_1), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2092_1_i) );
// C_///AND/D      x108y91     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2093_4 ( .OUT(na2093_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2093_5 ( .OUT(na2093_2), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2093_2_i) );
// C_AND/D///      x106y71     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2094_1 ( .OUT(na2094_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2094_2 ( .OUT(na2094_1), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2094_1_i) );
// C_///AND/D      x103y65     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2095_4 ( .OUT(na2095_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2095_5 ( .OUT(na2095_2), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2095_2_i) );
// C_AND/D///      x86y72     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2096_1 ( .OUT(na2096_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2096_2 ( .OUT(na2096_1), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2096_1_i) );
// C_///AND/D      x94y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2097_4 ( .OUT(na2097_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2097_5 ( .OUT(na2097_2), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2097_2_i) );
// C_AND/D///      x93y62     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2098_1 ( .OUT(na2098_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2098_2 ( .OUT(na2098_1), .CLK(1'b0), .EN(na1421_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2098_1_i) );
// C_///AND/D      x120y83     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2099_4 ( .OUT(na2099_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2099_5 ( .OUT(na2099_2), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2099_2_i) );
// C_AND/D///      x132y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2100_1 ( .OUT(na2100_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2100_2 ( .OUT(na2100_1), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2100_1_i) );
// C_///AND/D      x114y93     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2101_4 ( .OUT(na2101_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2101_5 ( .OUT(na2101_2), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2101_2_i) );
// C_AND/D///      x127y72     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2102_1 ( .OUT(na2102_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2102_2 ( .OUT(na2102_1), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2102_1_i) );
// C_///AND/D      x117y70     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2103_4 ( .OUT(na2103_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2103_5 ( .OUT(na2103_2), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2103_2_i) );
// C_AND/D///      x100y71     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2104_1 ( .OUT(na2104_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2104_2 ( .OUT(na2104_1), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2104_1_i) );
// C_///AND/D      x111y59     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2105_4 ( .OUT(na2105_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2105_5 ( .OUT(na2105_2), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2105_2_i) );
// C_///AND/D      x105y61     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2106_4 ( .OUT(na2106_2_i), .IN1(1'b1), .IN2(na3180_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2106_5 ( .OUT(na2106_2), .CLK(1'b0), .EN(na1423_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2106_2_i) );
// C_///AND/D      x104y89     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2107_4 ( .OUT(na2107_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2107_5 ( .OUT(na2107_2), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2107_2_i) );
// C_AND/D///      x128y89     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2108_1 ( .OUT(na2108_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2108_2 ( .OUT(na2108_1), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2108_1_i) );
// C_///AND/D      x122y97     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2109_4 ( .OUT(na2109_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2109_5 ( .OUT(na2109_2), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2109_2_i) );
// C_AND/D///      x116y71     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2110_1 ( .OUT(na2110_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2110_2 ( .OUT(na2110_1), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2110_1_i) );
// C_///AND/D      x112y71     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2111_4 ( .OUT(na2111_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2111_5 ( .OUT(na2111_2), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2111_2_i) );
// C_AND/D///      x87y80     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2112_1 ( .OUT(na2112_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2112_2 ( .OUT(na2112_1), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2112_1_i) );
// C_///AND/D      x114y65     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2113_4 ( .OUT(na2113_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2113_5 ( .OUT(na2113_2), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2113_2_i) );
// C_AND/D///      x109y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2114_1 ( .OUT(na2114_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2114_2 ( .OUT(na2114_1), .CLK(1'b0), .EN(na1424_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2114_1_i) );
// C_///AND/D      x117y95     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2115_4 ( .OUT(na2115_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2115_5 ( .OUT(na2115_2), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2115_2_i) );
// C_AND/D///      x130y100     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2116_1 ( .OUT(na2116_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2116_2 ( .OUT(na2116_1), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2116_1_i) );
// C_///AND/D      x125y102     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2117_4 ( .OUT(na2117_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2117_5 ( .OUT(na2117_2), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2117_2_i) );
// C_AND/D///      x123y86     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2118_1 ( .OUT(na2118_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2118_2 ( .OUT(na2118_1), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2118_1_i) );
// C_///AND/D      x113y83     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2119_4 ( .OUT(na2119_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2119_5 ( .OUT(na2119_2), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2119_2_i) );
// C_AND/D///      x99y84     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2120_1 ( .OUT(na2120_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2120_2 ( .OUT(na2120_1), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2120_1_i) );
// C_///AND/D      x105y58     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2121_4 ( .OUT(na2121_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2121_5 ( .OUT(na2121_2), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2121_2_i) );
// C_AND/D///      x117y62     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2122_1 ( .OUT(na2122_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2122_2 ( .OUT(na2122_1), .CLK(1'b0), .EN(na1426_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2122_1_i) );
// C_///AND/D      x97y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2123_4 ( .OUT(na2123_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2123_5 ( .OUT(na2123_2), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2123_2_i) );
// C_AND/D///      x120y92     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2124_1 ( .OUT(na2124_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2124_2 ( .OUT(na2124_1), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2124_1_i) );
// C_///AND/D      x119y97     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2125_4 ( .OUT(na2125_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2125_5 ( .OUT(na2125_2), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2125_2_i) );
// C_AND/D///      x110y72     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2126_1 ( .OUT(na2126_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2126_2 ( .OUT(na2126_1), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2126_1_i) );
// C_///AND/D      x101y68     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2127_4 ( .OUT(na2127_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2127_5 ( .OUT(na2127_2), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2127_2_i) );
// C_AND/D///      x85y71     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2128_1 ( .OUT(na2128_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2128_2 ( .OUT(na2128_1), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2128_1_i) );
// C_///AND/D      x98y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2129_4 ( .OUT(na2129_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2129_5 ( .OUT(na2129_2), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2129_2_i) );
// C_AND/D///      x103y60     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2130_1 ( .OUT(na2130_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2130_2 ( .OUT(na2130_1), .CLK(1'b0), .EN(na1427_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2130_1_i) );
// C_///AND/D      x93y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2131_4 ( .OUT(na2131_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2131_5 ( .OUT(na2131_2), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2131_2_i) );
// C_AND/D///      x113y93     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2132_1 ( .OUT(na2132_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2132_2 ( .OUT(na2132_1), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2132_1_i) );
// C_///AND/D      x113y93     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2133_4 ( .OUT(na2133_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2133_5 ( .OUT(na2133_2), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2133_2_i) );
// C_AND/D///      x107y75     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2134_1 ( .OUT(na2134_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2134_2 ( .OUT(na2134_1), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2134_1_i) );
// C_///AND/D      x91y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2135_4 ( .OUT(na2135_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2135_5 ( .OUT(na2135_2), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2135_2_i) );
// C_AND/D///      x81y78     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2136_1 ( .OUT(na2136_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2136_2 ( .OUT(na2136_1), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2136_1_i) );
// C_///AND/D      x93y58     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2137_4 ( .OUT(na2137_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2137_5 ( .OUT(na2137_2), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2137_2_i) );
// C_AND/D///      x95y60     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2138_1 ( .OUT(na2138_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2138_2 ( .OUT(na2138_1), .CLK(1'b0), .EN(na1428_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2138_1_i) );
// C_///AND/D      x118y94     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2139_4 ( .OUT(na2139_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2139_5 ( .OUT(na2139_2), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2139_2_i) );
// C_AND/D///      x131y100     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2140_1 ( .OUT(na2140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2140_2 ( .OUT(na2140_1), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2140_1_i) );
// C_///AND/D      x126y102     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2141_4 ( .OUT(na2141_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2141_5 ( .OUT(na2141_2), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2141_2_i) );
// C_AND/D///      x121y81     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2142_1 ( .OUT(na2142_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2142_2 ( .OUT(na2142_1), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2142_1_i) );
// C_///AND/D      x111y80     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2143_4 ( .OUT(na2143_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2143_5 ( .OUT(na2143_2), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2143_2_i) );
// C_AND/D///      x97y83     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2144_1 ( .OUT(na2144_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2144_2 ( .OUT(na2144_1), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2144_1_i) );
// C_///AND/D      x117y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2145_4 ( .OUT(na2145_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2145_5 ( .OUT(na2145_2), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2145_2_i) );
// C_AND/D///      x115y58     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2146_1 ( .OUT(na2146_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2146_2 ( .OUT(na2146_1), .CLK(1'b0), .EN(na1429_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2146_1_i) );
// C_///AND/D      x103y92     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2147_4 ( .OUT(na2147_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2147_5 ( .OUT(na2147_2), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2147_2_i) );
// C_AND/D///      x124y96     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2148_1 ( .OUT(na2148_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2148_2 ( .OUT(na2148_1), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2148_1_i) );
// C_///AND/D      x121y100     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2149_4 ( .OUT(na2149_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2149_5 ( .OUT(na2149_2), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2149_2_i) );
// C_AND/D///      x105y84     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2150_1 ( .OUT(na2150_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2150_2 ( .OUT(na2150_1), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2150_1_i) );
// C_///AND/D      x97y84     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2151_4 ( .OUT(na2151_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2151_5 ( .OUT(na2151_2), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2151_2_i) );
// C_AND/D///      x83y80     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2152_1 ( .OUT(na2152_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2152_2 ( .OUT(na2152_1), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2152_1_i) );
// C_///AND/D      x97y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2153_4 ( .OUT(na2153_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2153_5 ( .OUT(na2153_2), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2153_2_i) );
// C_AND/D///      x95y62     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2154_1 ( .OUT(na2154_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2154_2 ( .OUT(na2154_1), .CLK(1'b0), .EN(na1430_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2154_1_i) );
// C_///AND/D      x89y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2155_4 ( .OUT(na2155_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2155_5 ( .OUT(na2155_2), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2155_2_i) );
// C_AND/D///      x117y91     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2156_1 ( .OUT(na2156_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2156_2 ( .OUT(na2156_1), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2156_1_i) );
// C_///AND/D      x121y92     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2157_4 ( .OUT(na2157_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2157_5 ( .OUT(na2157_2), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2157_2_i) );
// C_AND/D///      x111y69     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2158_1 ( .OUT(na2158_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2158_2 ( .OUT(na2158_1), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2158_1_i) );
// C_///AND/D      x92y72     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2159_4 ( .OUT(na2159_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2159_5 ( .OUT(na2159_2), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2159_2_i) );
// C_AND/D///      x83y70     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2160_1 ( .OUT(na2160_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2160_2 ( .OUT(na2160_1), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2160_1_i) );
// C_///AND/D      x96y59     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2161_4 ( .OUT(na2161_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2161_5 ( .OUT(na2161_2), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2161_2_i) );
// C_AND/D///      x96y60     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2162_1 ( .OUT(na2162_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2162_2 ( .OUT(na2162_1), .CLK(1'b0), .EN(na1431_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2162_1_i) );
// C_///AND/D      x89y93     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2163_4 ( .OUT(na2163_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2163_5 ( .OUT(na2163_2), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2163_2_i) );
// C_AND/D///      x113y98     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2164_1 ( .OUT(na2164_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2164_2 ( .OUT(na2164_1), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2164_1_i) );
// C_///AND/D      x107y96     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2165_4 ( .OUT(na2165_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2165_5 ( .OUT(na2165_2), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2165_2_i) );
// C_AND/D///      x104y76     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2166_1 ( .OUT(na2166_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2166_2 ( .OUT(na2166_1), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2166_1_i) );
// C_AND/D///      x95y81     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2167_1 ( .OUT(na2167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3177_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2167_2 ( .OUT(na2167_1), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2167_1_i) );
// C_AND/D///      x81y75     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2168_1 ( .OUT(na2168_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2168_2 ( .OUT(na2168_1), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2168_1_i) );
// C_///AND/D      x89y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2169_4 ( .OUT(na2169_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2169_5 ( .OUT(na2169_2), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2169_2_i) );
// C_AND/D///      x92y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2170_1 ( .OUT(na2170_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2170_2 ( .OUT(na2170_1), .CLK(1'b0), .EN(na1432_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2170_1_i) );
// C_///AND/D      x101y90     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2171_4 ( .OUT(na2171_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2171_5 ( .OUT(na2171_2), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2171_2_i) );
// C_AND/D///      x118y96     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2172_1 ( .OUT(na2172_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2172_2 ( .OUT(na2172_1), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2172_1_i) );
// C_///AND/D      x122y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2173_4 ( .OUT(na2173_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2173_5 ( .OUT(na2173_2), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2173_2_i) );
// C_AND/D///      x109y84     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2174_1 ( .OUT(na2174_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2174_2 ( .OUT(na2174_1), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2174_1_i) );
// C_///AND/D      x99y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2175_4 ( .OUT(na2175_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2175_5 ( .OUT(na2175_2), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2175_2_i) );
// C_AND/D///      x89y82     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2176_1 ( .OUT(na2176_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2176_2 ( .OUT(na2176_1), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2176_1_i) );
// C_///AND/D      x99y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2177_4 ( .OUT(na2177_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2177_5 ( .OUT(na2177_2), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2177_2_i) );
// C_AND/D///      x99y66     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2178_1 ( .OUT(na2178_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2178_2 ( .OUT(na2178_1), .CLK(1'b0), .EN(na1433_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2178_1_i) );
// C_///AND/D      x91y86     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2179_4 ( .OUT(na2179_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2179_5 ( .OUT(na2179_2), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2179_2_i) );
// C_AND/D///      x115y95     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2180_1 ( .OUT(na2180_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2180_2 ( .OUT(na2180_1), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2180_1_i) );
// C_///AND/D      x107y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2181_4 ( .OUT(na2181_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2181_5 ( .OUT(na2181_2), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2181_2_i) );
// C_AND/D///      x109y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2182_1 ( .OUT(na2182_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2182_2 ( .OUT(na2182_1), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2182_1_i) );
// C_///AND/D      x95y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2183_4 ( .OUT(na2183_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2183_5 ( .OUT(na2183_2), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2183_2_i) );
// C_AND/D///      x85y77     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2184_1 ( .OUT(na2184_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2184_2 ( .OUT(na2184_1), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2184_1_i) );
// C_///AND/D      x96y62     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2185_4 ( .OUT(na2185_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2185_5 ( .OUT(na2185_2), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2185_2_i) );
// C_AND/D///      x93y60     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2186_1 ( .OUT(na2186_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2186_2 ( .OUT(na2186_1), .CLK(1'b0), .EN(na1434_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2186_1_i) );
// C_///AND/D      x118y95     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2187_4 ( .OUT(na2187_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2187_5 ( .OUT(na2187_2), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2187_2_i) );
// C_AND/D///      x122y104     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2188_1 ( .OUT(na2188_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2188_2 ( .OUT(na2188_1), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2188_1_i) );
// C_///AND/D      x129y104     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2189_4 ( .OUT(na2189_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2189_5 ( .OUT(na2189_2), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2189_2_i) );
// C_AND/D///      x121y86     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2190_1 ( .OUT(na2190_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2190_2 ( .OUT(na2190_1), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2190_1_i) );
// C_///AND/D      x115y80     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2191_4 ( .OUT(na2191_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2191_5 ( .OUT(na2191_2), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2191_2_i) );
// C_AND/D///      x99y78     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2192_1 ( .OUT(na2192_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2192_2 ( .OUT(na2192_1), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2192_1_i) );
// C_///AND/D      x106y62     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2193_4 ( .OUT(na2193_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2193_5 ( .OUT(na2193_2), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2193_2_i) );
// C_AND/D///      x114y61     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2194_1 ( .OUT(na2194_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2194_2 ( .OUT(na2194_1), .CLK(1'b0), .EN(na1435_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2194_1_i) );
// C_///AND/D      x103y93     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2195_4 ( .OUT(na2195_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2195_5 ( .OUT(na2195_2), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2195_2_i) );
// C_AND/D///      x127y92     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2196_1 ( .OUT(na2196_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2196_2 ( .OUT(na2196_1), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2196_1_i) );
// C_///AND/D      x121y97     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2197_4 ( .OUT(na2197_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2197_5 ( .OUT(na2197_2), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2197_2_i) );
// C_AND/D///      x111y84     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2198_1 ( .OUT(na2198_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2198_2 ( .OUT(na2198_1), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2198_1_i) );
// C_///AND/D      x98y86     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2199_4 ( .OUT(na2199_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2199_5 ( .OUT(na2199_2), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2199_2_i) );
// C_AND/D///      x89y81     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2200_1 ( .OUT(na2200_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2200_2 ( .OUT(na2200_1), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2200_1_i) );
// C_///AND/D      x106y64     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2201_4 ( .OUT(na2201_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2201_5 ( .OUT(na2201_2), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2201_2_i) );
// C_AND/D///      x103y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2202_1 ( .OUT(na2202_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2202_2 ( .OUT(na2202_1), .CLK(1'b0), .EN(na1436_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2202_1_i) );
// C_///AND/D      x93y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2203_4 ( .OUT(na2203_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2203_5 ( .OUT(na2203_2), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2203_2_i) );
// C_AND/D///      x113y92     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2204_1 ( .OUT(na2204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2204_2 ( .OUT(na2204_1), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2204_1_i) );
// C_///AND/D      x118y91     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2205_4 ( .OUT(na2205_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2205_5 ( .OUT(na2205_2), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2205_2_i) );
// C_AND/D///      x109y72     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2206_1 ( .OUT(na2206_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2206_2 ( .OUT(na2206_1), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2206_1_i) );
// C_///AND/D      x101y74     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2207_4 ( .OUT(na2207_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2207_5 ( .OUT(na2207_2), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2207_2_i) );
// C_AND/D///      x85y78     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2208_1 ( .OUT(na2208_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2208_2 ( .OUT(na2208_1), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2208_1_i) );
// C_///AND/D      x99y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2209_4 ( .OUT(na2209_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2209_5 ( .OUT(na2209_2), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2209_2_i) );
// C_AND/D///      x98y62     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2210_1 ( .OUT(na2210_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2210_2 ( .OUT(na2210_1), .CLK(1'b0), .EN(na1437_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2210_1_i) );
// C_///AND/D      x93y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2211_4 ( .OUT(na2211_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2211_5 ( .OUT(na2211_2), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2211_2_i) );
// C_AND/D///      x121y90     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2212_1 ( .OUT(na2212_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2212_2 ( .OUT(na2212_1), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2212_1_i) );
// C_///AND/D      x111y93     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2213_4 ( .OUT(na2213_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2213_5 ( .OUT(na2213_2), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2213_2_i) );
// C_AND/D///      x111y74     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2214_1 ( .OUT(na2214_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2214_2 ( .OUT(na2214_1), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2214_1_i) );
// C_///AND/D      x94y77     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2215_4 ( .OUT(na2215_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2215_5 ( .OUT(na2215_2), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2215_2_i) );
// C_AND/D///      x87y78     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2216_1 ( .OUT(na2216_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2216_2 ( .OUT(na2216_1), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2216_1_i) );
// C_///AND/D      x96y64     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2217_4 ( .OUT(na2217_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2217_5 ( .OUT(na2217_2), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2217_2_i) );
// C_AND/D///      x95y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2218_1 ( .OUT(na2218_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2218_2 ( .OUT(na2218_1), .CLK(1'b0), .EN(na1438_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2218_1_i) );
// C_///AND/D      x113y91     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2219_4 ( .OUT(na2219_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2219_5 ( .OUT(na2219_2), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2219_2_i) );
// C_AND/D///      x121y99     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2220_1 ( .OUT(na2220_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2220_2 ( .OUT(na2220_1), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2220_1_i) );
// C_///AND/D      x123y102     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2221_4 ( .OUT(na2221_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2221_5 ( .OUT(na2221_2), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2221_2_i) );
// C_AND/D///      x122y82     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2222_1 ( .OUT(na2222_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2222_2 ( .OUT(na2222_1), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2222_1_i) );
// C_///AND/D      x111y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2223_4 ( .OUT(na2223_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2223_5 ( .OUT(na2223_2), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2223_2_i) );
// C_AND/D///      x95y85     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2224_1 ( .OUT(na2224_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2224_2 ( .OUT(na2224_1), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2224_1_i) );
// C_///AND/D      x108y64     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2225_4 ( .OUT(na2225_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2225_5 ( .OUT(na2225_2), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2225_2_i) );
// C_AND/D///      x109y63     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2226_1 ( .OUT(na2226_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2226_2 ( .OUT(na2226_1), .CLK(1'b0), .EN(na1439_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2226_1_i) );
// C_///AND/D      x96y86     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2227_4 ( .OUT(na2227_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2227_5 ( .OUT(na2227_2), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2227_2_i) );
// C_///AND/D      x117y98     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2228_4 ( .OUT(na2228_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2228_5 ( .OUT(na2228_2), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2228_2_i) );
// C_///AND/D      x121y93     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2229_4 ( .OUT(na2229_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2229_5 ( .OUT(na2229_2), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2229_2_i) );
// C_AND/D///      x114y69     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2230_1 ( .OUT(na2230_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2230_2 ( .OUT(na2230_1), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2230_1_i) );
// C_///AND/D      x93y72     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2231_4 ( .OUT(na2231_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2231_5 ( .OUT(na2231_2), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2231_2_i) );
// C_AND/D///      x80y72     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2232_1 ( .OUT(na2232_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2232_2 ( .OUT(na2232_1), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2232_1_i) );
// C_///AND/D      x97y59     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2233_4 ( .OUT(na2233_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2233_5 ( .OUT(na2233_2), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2233_2_i) );
// C_AND/D///      x97y58     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2234_1 ( .OUT(na2234_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2234_2 ( .OUT(na2234_1), .CLK(1'b0), .EN(na1440_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2234_1_i) );
// C_///AND/D      x112y96     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2235_4 ( .OUT(na2235_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2235_5 ( .OUT(na2235_2), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2235_2_i) );
// C_AND/D///      x127y102     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2236_1 ( .OUT(na2236_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2236_2 ( .OUT(na2236_1), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2236_1_i) );
// C_///AND/D      x129y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2237_4 ( .OUT(na2237_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2237_5 ( .OUT(na2237_2), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2237_2_i) );
// C_AND/D///      x122y85     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2238_1 ( .OUT(na2238_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2238_2 ( .OUT(na2238_1), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2238_1_i) );
// C_///AND/D      x111y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2239_4 ( .OUT(na2239_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2239_5 ( .OUT(na2239_2), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2239_2_i) );
// C_AND/D///      x95y82     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2240_1 ( .OUT(na2240_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2240_2 ( .OUT(na2240_1), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2240_1_i) );
// C_///AND/D      x103y59     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2241_4 ( .OUT(na2241_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2241_5 ( .OUT(na2241_2), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2241_2_i) );
// C_AND/D///      x113y59     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2242_1 ( .OUT(na2242_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2242_2 ( .OUT(na2242_1), .CLK(1'b0), .EN(na1441_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2242_1_i) );
// C_///AND/D      x107y94     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2243_4 ( .OUT(na2243_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2243_5 ( .OUT(na2243_2), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2243_2_i) );
// C_AND/D///      x120y97     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2244_1 ( .OUT(na2244_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2244_2 ( .OUT(na2244_1), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2244_1_i) );
// C_///AND/D      x122y101     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2245_4 ( .OUT(na2245_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2245_5 ( .OUT(na2245_2), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2245_2_i) );
// C_AND/D///      x106y82     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2246_1 ( .OUT(na2246_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2246_2 ( .OUT(na2246_1), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2246_1_i) );
// C_///AND/D      x97y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2247_4 ( .OUT(na2247_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2247_5 ( .OUT(na2247_2), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2247_2_i) );
// C_AND/D///      x85y84     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2248_1 ( .OUT(na2248_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2248_2 ( .OUT(na2248_1), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2248_1_i) );
// C_///AND/D      x101y62     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2249_4 ( .OUT(na2249_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2249_5 ( .OUT(na2249_2), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2249_2_i) );
// C_AND/D///      x95y63     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2250_1 ( .OUT(na2250_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2250_2 ( .OUT(na2250_1), .CLK(1'b0), .EN(na1442_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2250_1_i) );
// C_///AND/D      x95y80     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2251_4 ( .OUT(na2251_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2251_5 ( .OUT(na2251_2), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2251_2_i) );
// C_AND/D///      x119y94     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2252_1 ( .OUT(na2252_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2252_2 ( .OUT(na2252_1), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2252_1_i) );
// C_///AND/D      x123y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2253_4 ( .OUT(na2253_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2253_5 ( .OUT(na2253_2), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2253_2_i) );
// C_AND/D///      x111y72     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2254_1 ( .OUT(na2254_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2254_2 ( .OUT(na2254_1), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2254_1_i) );
// C_///AND/D      x93y71     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2255_4 ( .OUT(na2255_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2255_5 ( .OUT(na2255_2), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2255_2_i) );
// C_AND/D///      x79y70     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2256_1 ( .OUT(na2256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2256_2 ( .OUT(na2256_1), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2256_1_i) );
// C_///AND/D      x91y58     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2257_4 ( .OUT(na2257_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2257_5 ( .OUT(na2257_2), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2257_2_i) );
// C_AND/D///      x95y58     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2258_1 ( .OUT(na2258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2258_2 ( .OUT(na2258_1), .CLK(1'b0), .EN(na1443_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2258_1_i) );
// C_///AND/D      x91y88     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2259_4 ( .OUT(na2259_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2259_5 ( .OUT(na2259_2), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2259_2_i) );
// C_AND/D///      x113y96     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2260_1 ( .OUT(na2260_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2260_2 ( .OUT(na2260_1), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2260_1_i) );
// C_///AND/D      x111y95     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2261_4 ( .OUT(na2261_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2261_5 ( .OUT(na2261_2), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2261_2_i) );
// C_AND/D///      x107y77     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2262_1 ( .OUT(na2262_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2262_2 ( .OUT(na2262_1), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2262_1_i) );
// C_///AND/D      x93y80     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2263_4 ( .OUT(na2263_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2263_5 ( .OUT(na2263_2), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2263_2_i) );
// C_AND/D///      x83y77     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2264_1 ( .OUT(na2264_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2264_2 ( .OUT(na2264_1), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2264_1_i) );
// C_///AND/D      x91y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2265_4 ( .OUT(na2265_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2265_5 ( .OUT(na2265_2), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2265_2_i) );
// C_AND/D///      x91y60     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2266_1 ( .OUT(na2266_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2266_2 ( .OUT(na2266_1), .CLK(1'b0), .EN(na1444_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2266_1_i) );
// C_///AND/D      x112y98     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2267_4 ( .OUT(na2267_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2267_5 ( .OUT(na2267_2), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2267_2_i) );
// C_AND/D///      x123y101     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2268_1 ( .OUT(na2268_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2268_2 ( .OUT(na2268_1), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2268_1_i) );
// C_///AND/D      x127y104     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2269_4 ( .OUT(na2269_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2269_5 ( .OUT(na2269_2), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2269_2_i) );
// C_AND/D///      x116y88     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2270_1 ( .OUT(na2270_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2270_2 ( .OUT(na2270_1), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2270_1_i) );
// C_///AND/D      x119y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2271_4 ( .OUT(na2271_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2271_5 ( .OUT(na2271_2), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2271_2_i) );
// C_AND/D///      x92y84     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2272_1 ( .OUT(na2272_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2272_2 ( .OUT(na2272_1), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2272_1_i) );
// C_///AND/D      x101y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2273_4 ( .OUT(na2273_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2273_5 ( .OUT(na2273_2), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2273_2_i) );
// C_AND/D///      x113y61     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2274_1 ( .OUT(na2274_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2274_2 ( .OUT(na2274_1), .CLK(1'b0), .EN(na1445_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2274_1_i) );
// C_///AND/D      x101y97     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2275_4 ( .OUT(na2275_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2275_5 ( .OUT(na2275_2), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2275_2_i) );
// C_AND/D///      x123y100     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2276_1 ( .OUT(na2276_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2276_2 ( .OUT(na2276_1), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2276_1_i) );
// C_///AND/D      x123y103     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2277_4 ( .OUT(na2277_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2277_5 ( .OUT(na2277_2), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2277_2_i) );
// C_AND/D///      x101y82     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2278_1 ( .OUT(na2278_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2278_2 ( .OUT(na2278_1), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2278_1_i) );
// C_///AND/D      x97y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2279_4 ( .OUT(na2279_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2279_5 ( .OUT(na2279_2), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2279_2_i) );
// C_AND/D///      x89y83     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2280_1 ( .OUT(na2280_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2280_2 ( .OUT(na2280_1), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2280_1_i) );
// C_///AND/D      x101y64     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2281_4 ( .OUT(na2281_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2281_5 ( .OUT(na2281_2), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2281_2_i) );
// C_AND/D///      x95y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2282_1 ( .OUT(na2282_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2282_2 ( .OUT(na2282_1), .CLK(1'b0), .EN(na1446_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2282_1_i) );
// C_///AND/D      x93y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2283_4 ( .OUT(na2283_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2283_5 ( .OUT(na2283_2), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2283_2_i) );
// C_AND/D///      x121y94     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2284_1 ( .OUT(na2284_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2284_2 ( .OUT(na2284_1), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2284_1_i) );
// C_///AND/D      x114y98     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2285_4 ( .OUT(na2285_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2285_5 ( .OUT(na2285_2), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2285_2_i) );
// C_AND/D///      x103y80     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2286_1 ( .OUT(na2286_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2286_2 ( .OUT(na2286_1), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2286_1_i) );
// C_///AND/D      x93y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2287_4 ( .OUT(na2287_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2287_5 ( .OUT(na2287_2), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2287_2_i) );
// C_AND/D///      x84y76     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2288_1 ( .OUT(na2288_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2288_2 ( .OUT(na2288_1), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2288_1_i) );
// C_AND/D///      x91y61     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2289_1 ( .OUT(na2289_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3179_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2289_2 ( .OUT(na2289_1), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2289_1_i) );
// C_AND/D///      x97y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2290_1 ( .OUT(na2290_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2290_2 ( .OUT(na2290_1), .CLK(1'b0), .EN(na1447_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2290_1_i) );
// C_///AND/D      x102y68     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2355_4 ( .OUT(na2355_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na214_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2355_5 ( .OUT(na2355_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2355_2_i) );
// C_AND/D///      x117y69     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2356_1 ( .OUT(na2356_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na264_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2356_2 ( .OUT(na2356_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2356_1_i) );
// C_///AND/D      x126y74     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2357_4 ( .OUT(na2357_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na277_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2357_5 ( .OUT(na2357_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2357_2_i) );
// C_AND/D///      x120y61     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2358_1 ( .OUT(na2358_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na287_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2358_2 ( .OUT(na2358_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2358_1_i) );
// C_///AND/D      x101y66     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2359_4 ( .OUT(na2359_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na295_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2359_5 ( .OUT(na2359_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2359_2_i) );
// C_AND/D///      x122y59     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2360_1 ( .OUT(na2360_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na300_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2360_2 ( .OUT(na2360_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2360_1_i) );
// C_///AND/D      x137y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2361_4 ( .OUT(na2361_2_i), .IN1(1'b1), .IN2(na309_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2361_5 ( .OUT(na2361_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2361_2_i) );
// C_AND/D///      x116y60     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2362_1 ( .OUT(na2362_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na315_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2362_2 ( .OUT(na2362_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2362_1_i) );
// C_///AND/D      x139y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2363_4 ( .OUT(na2363_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na972_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2363_5 ( .OUT(na2363_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2363_2_i) );
// C_AND/D///      x140y92     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2364_1 ( .OUT(na2364_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1018_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2364_2 ( .OUT(na2364_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2364_1_i) );
// C_///AND/D      x143y95     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2365_4 ( .OUT(na2365_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1030_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2365_5 ( .OUT(na2365_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2365_2_i) );
// C_AND/D///      x141y92     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2366_1 ( .OUT(na2366_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1035_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2366_2 ( .OUT(na2366_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2366_1_i) );
// C_///AND/D      x129y86     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2367_4 ( .OUT(na2367_2_i), .IN1(na1041_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2367_5 ( .OUT(na2367_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2367_2_i) );
// C_AND/D///      x133y89     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2368_1 ( .OUT(na2368_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1045_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2368_2 ( .OUT(na2368_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2368_1_i) );
// C_///AND/D      x138y71     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2369_4 ( .OUT(na2369_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1049_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2369_5 ( .OUT(na2369_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2369_2_i) );
// C_AND/D///      x135y78     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2370_1 ( .OUT(na2370_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1051_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2370_2 ( .OUT(na2370_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2370_1_i) );
// C_///AND/D      x140y98     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2371_4 ( .OUT(na2371_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na895_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2371_5 ( .OUT(na2371_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2371_2_i) );
// C_AND/D///      x135y98     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2372_1 ( .OUT(na2372_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4285_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2372_2 ( .OUT(na2372_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2372_1_i) );
// C_///AND/D      x152y93     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2373_4 ( .OUT(na2373_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na949_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2373_5 ( .OUT(na2373_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2373_2_i) );
// C_AND/D///      x152y95     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2374_1 ( .OUT(na2374_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na955_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2374_2 ( .OUT(na2374_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2374_1_i) );
// C_///AND/D      x146y96     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2375_4 ( .OUT(na2375_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na962_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2375_5 ( .OUT(na2375_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2375_2_i) );
// C_AND/D///      x146y94     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2376_1 ( .OUT(na2376_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na965_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2376_2 ( .OUT(na2376_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2376_1_i) );
// C_///AND/D      x143y88     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2377_4 ( .OUT(na2377_2_i), .IN1(1'b1), .IN2(na968_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2377_5 ( .OUT(na2377_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2377_2_i) );
// C_AND/D///      x145y80     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2378_1 ( .OUT(na2378_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na970_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2378_2 ( .OUT(na2378_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2378_1_i) );
// C_///AND/D      x124y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2379_4 ( .OUT(na2379_2_i), .IN1(1'b1), .IN2(na816_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2379_5 ( .OUT(na2379_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2379_2_i) );
// C_AND/D///      x112y82     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2380_1 ( .OUT(na2380_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na862_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2380_2 ( .OUT(na2380_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2380_1_i) );
// C_///AND/D      x124y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2381_4 ( .OUT(na2381_2_i), .IN1(1'b1), .IN2(na871_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2381_5 ( .OUT(na2381_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2381_2_i) );
// C_AND/D///      x129y76     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2382_1 ( .OUT(na2382_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na877_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2382_2 ( .OUT(na2382_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2382_1_i) );
// C_///AND/D      x111y71     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2383_4 ( .OUT(na2383_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2383_5 ( .OUT(na2383_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2383_2_i) );
// C_AND/D///      x120y70     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2384_1 ( .OUT(na2384_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na887_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2384_2 ( .OUT(na2384_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2384_1_i) );
// C_///AND/D      x126y68     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2385_4 ( .OUT(na2385_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2385_5 ( .OUT(na2385_2), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2385_2_i) );
// C_AND/D///      x126y66     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2386_1 ( .OUT(na2386_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na892_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2386_2 ( .OUT(na2386_1), .CLK(1'b0), .EN(na1450_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2386_1_i) );
// C_///AND/D      x124y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2402_4 ( .OUT(na2402_2_i), .IN1(1'b1), .IN2(na816_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2402_5 ( .OUT(na2402_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2402_2_i) );
// C_AND/D///      x110y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2403_1 ( .OUT(na2403_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na862_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2403_2 ( .OUT(na2403_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2403_1_i) );
// C_///AND/D      x129y84     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2404_4 ( .OUT(na2404_2_i), .IN1(1'b1), .IN2(na871_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2404_5 ( .OUT(na2404_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2404_2_i) );
// C_AND/D///      x138y70     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2405_1 ( .OUT(na2405_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na877_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2405_2 ( .OUT(na2405_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2405_1_i) );
// C_///AND/D      x114y76     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2406_4 ( .OUT(na2406_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2406_5 ( .OUT(na2406_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2406_2_i) );
// C_AND/D///      x129y70     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2407_1 ( .OUT(na2407_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na887_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2407_2 ( .OUT(na2407_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2407_1_i) );
// C_///AND/D      x137y66     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2408_4 ( .OUT(na2408_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2408_5 ( .OUT(na2408_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2408_2_i) );
// C_AND/D///      x135y65     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2409_1 ( .OUT(na2409_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na892_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2409_2 ( .OUT(na2409_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2409_1_i) );
// C_///AND/D      x114y74     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2410_4 ( .OUT(na2410_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na214_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2410_5 ( .OUT(na2410_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2410_2_i) );
// C_AND/D///      x125y75     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2411_1 ( .OUT(na2411_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na264_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2411_2 ( .OUT(na2411_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2411_1_i) );
// C_///AND/D      x128y77     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2412_4 ( .OUT(na2412_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na277_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2412_5 ( .OUT(na2412_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2412_2_i) );
// C_AND/D///      x122y61     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2413_1 ( .OUT(na2413_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na287_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2413_2 ( .OUT(na2413_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2413_1_i) );
// C_///AND/D      x116y66     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2414_4 ( .OUT(na2414_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na295_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2414_5 ( .OUT(na2414_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2414_2_i) );
// C_AND/D///      x125y66     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2415_1 ( .OUT(na2415_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na300_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2415_2 ( .OUT(na2415_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2415_1_i) );
// C_///AND/D      x141y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2416_4 ( .OUT(na2416_2_i), .IN1(1'b1), .IN2(na309_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2416_5 ( .OUT(na2416_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2416_2_i) );
// C_AND/D///      x116y62     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2417_1 ( .OUT(na2417_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na315_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2417_2 ( .OUT(na2417_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2417_1_i) );
// C_///AND/D      x133y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2418_4 ( .OUT(na2418_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na972_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2418_5 ( .OUT(na2418_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2418_2_i) );
// C_AND/D///      x142y91     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2419_1 ( .OUT(na2419_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1018_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2419_2 ( .OUT(na2419_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2419_1_i) );
// C_///AND/D      x134y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2420_4 ( .OUT(na2420_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1030_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2420_5 ( .OUT(na2420_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2420_2_i) );
// C_AND/D///      x135y91     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2421_1 ( .OUT(na2421_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1035_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2421_2 ( .OUT(na2421_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2421_1_i) );
// C_///AND/D      x127y83     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2422_4 ( .OUT(na2422_2_i), .IN1(na1041_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2422_5 ( .OUT(na2422_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2422_2_i) );
// C_AND/D///      x129y87     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2423_1 ( .OUT(na2423_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1045_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2423_2 ( .OUT(na2423_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2423_1_i) );
// C_///AND/D      x134y77     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2424_4 ( .OUT(na2424_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1049_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2424_5 ( .OUT(na2424_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2424_2_i) );
// C_AND/D///      x135y77     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2425_1 ( .OUT(na2425_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1051_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2425_2 ( .OUT(na2425_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2425_1_i) );
// C_///AND/D      x148y96     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2426_4 ( .OUT(na2426_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na895_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2426_5 ( .OUT(na2426_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2426_2_i) );
// C_AND/D///      x137y97     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2427_1 ( .OUT(na2427_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4285_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2427_2 ( .OUT(na2427_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2427_1_i) );
// C_///AND/D      x154y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2428_4 ( .OUT(na2428_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na949_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2428_5 ( .OUT(na2428_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2428_2_i) );
// C_///AND/D      x156y93     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2429_4 ( .OUT(na2429_2_i), .IN1(na955_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2429_5 ( .OUT(na2429_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2429_2_i) );
// C_///AND/D      x154y98     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2430_4 ( .OUT(na2430_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na962_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2430_5 ( .OUT(na2430_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2430_2_i) );
// C_AND/D///      x149y91     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2431_1 ( .OUT(na2431_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na965_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2431_2 ( .OUT(na2431_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2431_1_i) );
// C_///AND/D      x143y81     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2432_4 ( .OUT(na2432_2_i), .IN1(1'b1), .IN2(na968_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2432_5 ( .OUT(na2432_2), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2432_2_i) );
// C_AND/D///      x147y79     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2433_1 ( .OUT(na2433_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na970_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2433_2 ( .OUT(na2433_1), .CLK(1'b0), .EN(na349_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2433_1_i) );
// C_///AND/D      x140y72     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2918_4 ( .OUT(na2918_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1141_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2918_5 ( .OUT(na2918_2), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2918_2_i) );
// C_AND/D///      x142y74     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2919_1 ( .OUT(na2919_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1143_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2919_2 ( .OUT(na2919_1), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2919_1_i) );
// C_///AND/D      x145y77     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2920_4 ( .OUT(na2920_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1144_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2920_5 ( .OUT(na2920_2), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2920_2_i) );
// C_AND/D///      x140y68     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2921_1 ( .OUT(na2921_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2921_2 ( .OUT(na2921_1), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2921_1_i) );
// C_///AND/D      x140y68     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2922_4 ( .OUT(na2922_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1146_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2922_5 ( .OUT(na2922_2), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2922_2_i) );
// C_AND/D///      x135y72     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2923_1 ( .OUT(na2923_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1147_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2923_2 ( .OUT(na2923_1), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2923_1_i) );
// C_///AND/D      x143y67     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2924_4 ( .OUT(na2924_2_i), .IN1(1'b1), .IN2(na1148_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2924_5 ( .OUT(na2924_2), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2924_2_i) );
// C_AND/D///      x137y68     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2925_1 ( .OUT(na2925_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1149_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2925_2 ( .OUT(na2925_1), .CLK(1'b0), .EN(na26_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2925_1_i) );
// C_///AND/D      x132y92     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2926_4 ( .OUT(na2926_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na972_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2926_5 ( .OUT(na2926_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2926_2_i) );
// C_AND/D///      x145y91     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2927_1 ( .OUT(na2927_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1018_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2927_2 ( .OUT(na2927_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2927_1_i) );
// C_///AND/D      x148y94     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2928_4 ( .OUT(na2928_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1030_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2928_5 ( .OUT(na2928_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2928_2_i) );
// C_AND/D///      x145y93     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2929_1 ( .OUT(na2929_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1035_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2929_2 ( .OUT(na2929_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2929_1_i) );
// C_///AND/D      x138y92     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2930_4 ( .OUT(na2930_2_i), .IN1(na1041_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2930_5 ( .OUT(na2930_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2930_2_i) );
// C_AND/D///      x138y88     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2931_1 ( .OUT(na2931_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1045_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2931_2 ( .OUT(na2931_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2931_1_i) );
// C_///AND/D      x141y75     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2932_4 ( .OUT(na2932_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1049_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2932_5 ( .OUT(na2932_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2932_2_i) );
// C_AND/D///      x137y78     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2933_1 ( .OUT(na2933_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1051_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2933_2 ( .OUT(na2933_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2933_1_i) );
// C_///AND/D      x143y99     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2934_4 ( .OUT(na2934_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na895_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2934_5 ( .OUT(na2934_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2934_2_i) );
// C_AND/D///      x136y98     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2935_1 ( .OUT(na2935_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4285_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2935_2 ( .OUT(na2935_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2935_1_i) );
// C_///AND/D      x156y95     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2936_4 ( .OUT(na2936_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na949_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2936_5 ( .OUT(na2936_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2936_2_i) );
// C_AND/D///      x156y95     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2937_1 ( .OUT(na2937_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na955_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2937_2 ( .OUT(na2937_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2937_1_i) );
// C_///AND/D      x154y91     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2938_4 ( .OUT(na2938_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na962_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2938_5 ( .OUT(na2938_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2938_2_i) );
// C_AND/D///      x154y94     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2939_1 ( .OUT(na2939_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na965_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2939_2 ( .OUT(na2939_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2939_1_i) );
// C_///AND/D      x148y90     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2940_4 ( .OUT(na2940_2_i), .IN1(1'b1), .IN2(na968_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2940_5 ( .OUT(na2940_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2940_2_i) );
// C_AND/D///      x148y79     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2941_1 ( .OUT(na2941_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na970_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2941_2 ( .OUT(na2941_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2941_1_i) );
// C_///AND/D      x119y73     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2942_4 ( .OUT(na2942_2_i), .IN1(1'b1), .IN2(na816_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2942_5 ( .OUT(na2942_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2942_2_i) );
// C_AND/D///      x111y86     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2943_1 ( .OUT(na2943_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na862_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2943_2 ( .OUT(na2943_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2943_1_i) );
// C_///AND/D      x121y82     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2944_4 ( .OUT(na2944_2_i), .IN1(1'b1), .IN2(na871_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2944_5 ( .OUT(na2944_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2944_2_i) );
// C_AND/D///      x127y74     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2945_1 ( .OUT(na2945_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na877_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2945_2 ( .OUT(na2945_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2945_1_i) );
// C_///AND/D      x114y71     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2946_4 ( .OUT(na2946_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2946_5 ( .OUT(na2946_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2946_2_i) );
// C_AND/D///      x118y72     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2947_1 ( .OUT(na2947_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na887_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2947_2 ( .OUT(na2947_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2947_1_i) );
// C_///AND/D      x126y67     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2948_4 ( .OUT(na2948_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2948_5 ( .OUT(na2948_2), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2948_2_i) );
// C_AND/D///      x123y65     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2949_1 ( .OUT(na2949_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na892_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2949_2 ( .OUT(na2949_1), .CLK(1'b0), .EN(na1451_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2949_1_i) );
// C_///AND/D      x139y69     80'h40_EC00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3142_4 ( .OUT(na3142_2_i), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3142_5 ( .OUT(na3142_2), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3142_2_i) );
// C_AND/D///      x139y62     80'h40_EC00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3143_1 ( .OUT(na3143_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1335_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3143_2 ( .OUT(na3143_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3143_1_i) );
// C_///AND/D      x146y68     80'h40_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3144_4 ( .OUT(na3144_2_i), .IN1(na1335_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3144_5 ( .OUT(na3144_2), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3144_2_i) );
// C_AND/D///      x140y62     80'h40_EC00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3145_1 ( .OUT(na3145_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1336_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3145_2 ( .OUT(na3145_1), .CLK(1'b0), .EN(1'b1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3145_1_i) );
// C_///AND/D      x95y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3154_4 ( .OUT(na3154_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3154_5 ( .OUT(na3154_2), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3154_2_i) );
// C_AND/D///      x119y96     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3155_1 ( .OUT(na3155_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3155_2 ( .OUT(na3155_1), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3155_1_i) );
// C_///AND/D      x119y96     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3156_4 ( .OUT(na3156_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3156_5 ( .OUT(na3156_2), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3156_2_i) );
// C_AND/D///      x112y72     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3157_1 ( .OUT(na3157_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3157_2 ( .OUT(na3157_1), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3157_1_i) );
// C_///AND/D      x100y74     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3158_4 ( .OUT(na3158_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3158_5 ( .OUT(na3158_2), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3158_2_i) );
// C_AND/D///      x83y76     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3159_1 ( .OUT(na3159_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3159_2 ( .OUT(na3159_1), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3159_1_i) );
// C_///AND/D      x99y58     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3160_4 ( .OUT(na3160_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3160_5 ( .OUT(na3160_2), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3160_2_i) );
// C_AND/D///      x99y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3161_1 ( .OUT(na3161_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3161_2 ( .OUT(na3161_1), .CLK(1'b0), .EN(na1479_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3161_1_i) );
// C_///AND/D      x95y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3165_4 ( .OUT(na3165_2_i), .IN1(1'b1), .IN2(na3173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3165_5 ( .OUT(na3165_2), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3165_2_i) );
// C_AND/D///      x121y96     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3166_1 ( .OUT(na3166_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3174_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3166_2 ( .OUT(na3166_1), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3166_1_i) );
// C_///AND/D      x124y99     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3167_4 ( .OUT(na3167_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3175_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3167_5 ( .OUT(na3167_2), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3167_2_i) );
// C_AND/D///      x113y70     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3168_1 ( .OUT(na3168_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3168_2 ( .OUT(na3168_1), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3168_1_i) );
// C_///AND/D      x101y72     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3169_4 ( .OUT(na3169_2_i), .IN1(1'b1), .IN2(na3177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3169_5 ( .OUT(na3169_2), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3169_2_i) );
// C_AND/D///      x81y73     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3170_1 ( .OUT(na3170_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3170_2 ( .OUT(na3170_1), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3170_1_i) );
// C_///AND/D      x98y61     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3171_4 ( .OUT(na3171_2_i), .IN1(1'b1), .IN2(na3179_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3171_5 ( .OUT(na3171_2), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3171_2_i) );
// C_AND/D///      x101y58     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3172_1 ( .OUT(na3172_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3180_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3172_2 ( .OUT(na3172_1), .CLK(1'b0), .EN(na1477_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3172_1_i) );
// C_///AND/D      x107y92     80'h40_F800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3173_4 ( .OUT(na3173_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3173_5 ( .OUT(na3173_2), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3173_2_i) );
// C_AND/D///      x122y95     80'h40_F800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3174_1 ( .OUT(na3174_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3175_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3174_2 ( .OUT(na3174_1), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3174_1_i) );
// C_///AND/D      x122y95     80'h40_F800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3175_4 ( .OUT(na3175_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3176_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3175_5 ( .OUT(na3175_2), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3175_2_i) );
// C_AND/D///      x114y78     80'h40_F800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3176_1 ( .OUT(na3176_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3177_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3176_2 ( .OUT(na3176_1), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3176_1_i) );
// C_AND/D///      x107y78     80'h40_F800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3177_1 ( .OUT(na3177_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3177_2 ( .OUT(na3177_1), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3177_1_i) );
// C_AND/D///      x89y76     80'h40_F800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3178_1 ( .OUT(na3178_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3179_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3178_2 ( .OUT(na3178_1), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3178_1_i) );
// C_///AND/D      x105y60     80'h40_F800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3179_4 ( .OUT(na3179_2_i), .IN1(1'b1), .IN2(na3180_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3179_5 ( .OUT(na3179_2), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3179_2_i) );
// C_AND/D///      x97y60     80'h40_F800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3180_1 ( .OUT(na3180_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3223_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3180_2 ( .OUT(na3180_1), .CLK(1'b0), .EN(na1394_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3180_1_i) );
// C_///AND/D      x88y59     80'h40_E800_80_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3196_4 ( .OUT(na3196_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3196_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3196_5 ( .OUT(na3196_2), .CLK(1'b0), .EN(na1397_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3196_2_i) );
// C_AND/D///      x115y88     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3198_1 ( .OUT(na3198_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3173_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3198_2 ( .OUT(na3198_1), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3198_1_i) );
// C_///AND/D      x119y86     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3199_4 ( .OUT(na3199_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3199_5 ( .OUT(na3199_2), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3199_2_i) );
// C_AND/D///      x125y88     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3200_1 ( .OUT(na3200_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3175_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3200_2 ( .OUT(na3200_1), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3200_1_i) );
// C_///AND/D      x119y74     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3201_4 ( .OUT(na3201_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3176_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3201_5 ( .OUT(na3201_2), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3201_2_i) );
// C_AND/D///      x113y78     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3202_1 ( .OUT(na3202_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3177_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3202_2 ( .OUT(na3202_1), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3202_1_i) );
// C_///AND/D      x93y74     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3203_4 ( .OUT(na3203_2_i), .IN1(1'b1), .IN2(na3178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3203_5 ( .OUT(na3203_2), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3203_2_i) );
// C_AND/D///      x105y64     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3204_1 ( .OUT(na3204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3179_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3204_2 ( .OUT(na3204_1), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3204_1_i) );
// C_///AND/D      x119y60     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3205_4 ( .OUT(na3205_2_i), .IN1(1'b1), .IN2(na3180_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3205_5 ( .OUT(na3205_2), .CLK(1'b0), .EN(na1399_2), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3205_2_i) );
// C_AND/D///      x103y90     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3206_1 ( .OUT(na3206_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3173_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3206_2 ( .OUT(na3206_1), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3206_1_i) );
// C_///AND/D      x111y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3207_4 ( .OUT(na3207_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3207_5 ( .OUT(na3207_2), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3207_2_i) );
// C_AND/D///      x121y98     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3208_1 ( .OUT(na3208_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3175_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3208_2 ( .OUT(na3208_1), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3208_1_i) );
// C_///AND/D      x101y78     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3209_4 ( .OUT(na3209_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3176_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3209_5 ( .OUT(na3209_2), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3209_2_i) );
// C_AND/D///      x101y81     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3210_1 ( .OUT(na3210_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3177_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3210_2 ( .OUT(na3210_1), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3210_1_i) );
// C_///AND/D      x84y78     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3211_4 ( .OUT(na3211_2_i), .IN1(1'b1), .IN2(na3178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3211_5 ( .OUT(na3211_2), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3211_2_i) );
// C_AND/D///      x93y66     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3212_1 ( .OUT(na3212_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3179_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3212_2 ( .OUT(na3212_1), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3212_1_i) );
// C_///AND/D      x107y63     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3213_4 ( .OUT(na3213_2_i), .IN1(1'b1), .IN2(na3180_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3213_5 ( .OUT(na3213_2), .CLK(1'b0), .EN(na1478_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3213_2_i) );
// C_AND/D///      x85y59     80'h40_F800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3223_1 ( .OUT(na3223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3281_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3223_2 ( .OUT(na3223_1), .CLK(1'b0), .EN(na3289_1), .SR(1'b1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3223_1_i) );
// C_///AND/D      x153y61     80'h40_E800_80_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3235_4 ( .OUT(na3235_2_i), .IN1(~na3235_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3235_5 ( .OUT(na3235_2), .CLK(1'b0), .EN(na1391_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3235_2_i) );
// C_AND/D///      x104y88     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3237_1 ( .OUT(na3237_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3173_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3237_2 ( .OUT(na3237_1), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3237_1_i) );
// C_///AND/D      x109y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3238_4 ( .OUT(na3238_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3238_5 ( .OUT(na3238_2), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3238_2_i) );
// C_AND/D///      x127y98     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3239_1 ( .OUT(na3239_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3175_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3239_2 ( .OUT(na3239_1), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3239_1_i) );
// C_///AND/D      x102y80     80'h40_E800_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3240_4 ( .OUT(na3240_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3176_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3240_5 ( .OUT(na3240_2), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3240_2_i) );
// C_AND/D///      x102y80     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3241_1 ( .OUT(na3241_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3177_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3241_2 ( .OUT(na3241_1), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3241_1_i) );
// C_///AND/D      x81y76     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3242_4 ( .OUT(na3242_2_i), .IN1(1'b1), .IN2(na3178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3242_5 ( .OUT(na3242_2), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3242_2_i) );
// C_AND/D///      x100y67     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3243_1 ( .OUT(na3243_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3179_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a3243_2 ( .OUT(na3243_1), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3243_1_i) );
// C_///AND/D      x109y61     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3244_4 ( .OUT(na3244_2_i), .IN1(1'b1), .IN2(na3180_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a3244_5 ( .OUT(na3244_2), .CLK(1'b0), .EN(na1474_1), .SR(na3289_1), .CINY2(na4512_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3244_2_i) );
// C_MX2b////      x140y71     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3248_1 ( .OUT(na3248_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1819_1), .IN6(na1742_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x142y66     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3249_1 ( .OUT(na3249_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1744_2), .IN6(na1824_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x144y68     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3250_1 ( .OUT(na3250_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na279_1), .IN8(na1747_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x133y64     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3251_1 ( .OUT(na3251_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1829_1), .IN6(na1749_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x132y63     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3252_1 ( .OUT(na3252_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1751_1), .IN8(na1834_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x127y61     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3253_1 ( .OUT(na3253_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1838_1), .IN8(na1753_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y62     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3254_1 ( .OUT(na3254_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1755_1), .IN6(na1862_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y58     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3255_1 ( .OUT(na3255_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na316_1), .IN8(na1757_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x141y70     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3256_1 ( .OUT(na3256_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na324_1), .IN6(na1759_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x152y67     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3257_1 ( .OUT(na3257_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na333_1), .IN8(na1760_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x145y71     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3258_1 ( .OUT(na3258_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na342_1), .IN6(na1762_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y64     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3259_1 ( .OUT(na3259_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na353_1), .IN8(na1764_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y66     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3260_1 ( .OUT(na3260_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na362_1), .IN8(na1766_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x128y63     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3261_1 ( .OUT(na3261_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1768_1), .IN8(na371_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y61     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3262_1 ( .OUT(na3262_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1770_1), .IN8(na380_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y63     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3263_1 ( .OUT(na3263_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1772_1), .IN6(na389_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x148y72     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3264_1 ( .OUT(na3264_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1774_1), .IN8(na397_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x148y73     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3265_1 ( .OUT(na3265_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1775_1), .IN8(na405_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x150y71     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3266_1 ( .OUT(na3266_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1777_1), .IN6(na414_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x150y69     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3267_1 ( .OUT(na3267_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1779_1), .IN6(na423_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y67     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3268_1 ( .OUT(na3268_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1781_1), .IN6(na432_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x145y70     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3269_1 ( .OUT(na3269_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na441_1), .IN6(na1783_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x137y65     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3270_1 ( .OUT(na3270_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1784_1), .IN8(na449_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x144y64     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3271_1 ( .OUT(na3271_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na458_1), .IN8(na1785_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y72     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3272_1 ( .OUT(na3272_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na467_1), .IN8(na1787_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x146y71     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3273_1 ( .OUT(na3273_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na476_1), .IN6(na1789_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x147y71     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3274_1 ( .OUT(na3274_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1790_2), .IN8(na485_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x145y68     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3275_1 ( .OUT(na3275_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1791_1), .IN8(na494_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x142y68     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3276_1 ( .OUT(na3276_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na503_1), .IN6(na1793_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x143y65     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3277_1 ( .OUT(na3277_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1795_1), .IN6(na512_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y63     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3278_1 ( .OUT(na3278_1), .IN1(~na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1797_1), .IN6(na521_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x136y63     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3279_1 ( .OUT(na3279_1), .IN1(na1481_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na530_1), .IN6(na1798_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a3280 ( .Y(na3280_1), .I(clk) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a3281 ( .Y(na3281_1), .I(data_in) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3282 ( .O(data_out), .A(na4158_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3283 ( .O(led[0]), .A(na4159_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3284 ( .O(led[1]), .A(na4160_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3285 ( .O(led[2]), .A(na4161_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3286 ( .O(led[3]), .A(na4162_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3287 ( .O(led[4]), .A(na4163_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a3288 ( .O(led[5]), .A(na4164_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a3289 ( .Y(na3289_1), .I(reset_n) );
// C_AND///AND/      x106y81     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3290_1 ( .OUT(na3290_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(1'b1), .IN8(na776_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3290_4 ( .OUT(na3290_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na680_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y73     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3292_4 ( .OUT(na3292_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(na616_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y75     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3293_1 ( .OUT(na3293_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2083_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x115y75     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3294_4 ( .OUT(na3294_2), .IN1(~na1331_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1332_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x145y75     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3296_2 ( .OUT(na3296_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3296_6 ( .COUTY1(na3296_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3296_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x143y88     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3297_1 ( .OUT(na3297_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1870_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x126y81     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3298_1 ( .OUT(na3298_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(na681_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3298_4 ( .OUT(na3298_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na777_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y79     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3300_1 ( .OUT(na3300_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4350_2), .IN7(1'b1), .IN8(na2084_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y75     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3301_4 ( .OUT(na3301_2), .IN1(~na16_2), .IN2(1'b1), .IN3(na617_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x130y87     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3303_1 ( .OUT(na3303_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na778_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3303_4 ( .OUT(na3303_2), .IN1(na26_2), .IN2(na682_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y78     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3305_4 ( .OUT(na3305_2), .IN1(na618_1), .IN2(1'b1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y79     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3306_4 ( .OUT(na3306_2), .IN1(na16_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2085_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x132y74     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3308_1 ( .OUT(na3308_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na779_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3308_4 ( .OUT(na3308_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na683_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y65     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3310_1 ( .OUT(na3310_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na619_1), .IN7(na15_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x118y69     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3311_4 ( .OUT(na3311_2), .IN1(na16_2), .IN2(1'b1), .IN3(na2086_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x115y71     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3313_1 ( .OUT(na3313_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na780_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3313_4 ( .OUT(na3313_2), .IN1(na26_2), .IN2(na684_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y68     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3315_1 ( .OUT(na3315_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na15_2), .IN8(na620_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y67     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3316_4 ( .OUT(na3316_2), .IN1(na2087_2), .IN2(na4170_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x101y73     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3318_1 ( .OUT(na3318_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na781_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3318_4 ( .OUT(na3318_2), .IN1(na26_2), .IN2(1'b1), .IN3(na685_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y67     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3320_1 ( .OUT(na3320_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na621_1), .IN6(1'b1), .IN7(na15_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y71     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3321_1 ( .OUT(na3321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(na2088_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y65     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3323_1 ( .OUT(na3323_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(na686_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3323_4 ( .OUT(na3323_2), .IN1(na26_1), .IN2(na782_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x120y62     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3325_1 ( .OUT(na3325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2089_2), .IN7(1'b1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y67     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3326_4 ( .OUT(na3326_2), .IN1(~na16_2), .IN2(1'b1), .IN3(na622_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x112y68     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3328_1 ( .OUT(na3328_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na783_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3328_4 ( .OUT(na3328_2), .IN1(na26_2), .IN2(1'b1), .IN3(na687_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y63     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3330_1 ( .OUT(na3330_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na623_1), .IN7(na15_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y61     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3331_4 ( .OUT(na3331_2), .IN1(na2090_1), .IN2(na4170_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y82     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3333_1 ( .OUT(na3333_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(1'b1), .IN8(na784_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3333_4 ( .OUT(na3333_2), .IN1(na26_2), .IN2(1'b1), .IN3(na688_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y76     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3335_4 ( .OUT(na3335_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(na624_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y82     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3336_4 ( .OUT(na3336_2), .IN1(na2091_2), .IN2(na4170_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x126y86     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3338_1 ( .OUT(na3338_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na689_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3338_4 ( .OUT(na3338_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na785_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y78     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3340_4 ( .OUT(na3340_2), .IN1(na625_1), .IN2(1'b1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y82     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3341_1 ( .OUT(na3341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(na2092_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x118y88     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3343_1 ( .OUT(na3343_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na690_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3343_4 ( .OUT(na3343_2), .IN1(na26_1), .IN2(na786_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y79     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3345_4 ( .OUT(na3345_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(na626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y85     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3346_1 ( .OUT(na3346_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(na2093_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x109y76     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3348_1 ( .OUT(na3348_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(1'b1), .IN8(na787_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3348_4 ( .OUT(na3348_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na691_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y72     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3350_1 ( .OUT(na3350_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na627_1), .IN6(1'b1), .IN7(na15_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y71     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3351_1 ( .OUT(na3351_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(na2094_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x111y78     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3353_1 ( .OUT(na3353_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na692_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3353_4 ( .OUT(na3353_2), .IN1(na26_1), .IN2(1'b1), .IN3(na788_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x120y71     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3355_4 ( .OUT(na3355_2), .IN1(na2095_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y72     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3356_1 ( .OUT(na3356_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na16_2), .IN6(1'b1), .IN7(na628_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y76     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3358_1 ( .OUT(na3358_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(1'b1), .IN8(na789_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3358_4 ( .OUT(na3358_2), .IN1(na26_2), .IN2(na693_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y72     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3360_4 ( .OUT(na3360_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(na629_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y75     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3361_1 ( .OUT(na3361_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2096_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x104y70     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3363_1 ( .OUT(na3363_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(1'b1), .IN8(na790_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3363_4 ( .OUT(na3363_2), .IN1(na26_2), .IN2(na694_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y70     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3365_4 ( .OUT(na3365_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(na630_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y68     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3366_1 ( .OUT(na3366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(na2097_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x104y68     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3368_1 ( .OUT(na3368_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na791_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3368_4 ( .OUT(na3368_2), .IN1(na26_2), .IN2(na695_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y68     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3370_1 ( .OUT(na3370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na631_1), .IN7(na15_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y65     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3371_1 ( .OUT(na3371_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(na2098_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x135y93     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3373_1 ( .OUT(na3373_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na696_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3373_4 ( .OUT(na3373_2), .IN1(na26_1), .IN2(na792_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x132y88     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3375_4 ( .OUT(na3375_2), .IN1(1'b1), .IN2(na4350_2), .IN3(1'b1), .IN4(na1961_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y90     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3376_1 ( .OUT(na3376_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na632_1), .IN6(~na4170_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x133y93     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3378_1 ( .OUT(na3378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(1'b1), .IN8(na697_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3378_4 ( .OUT(na3378_2), .IN1(na26_1), .IN2(1'b1), .IN3(na793_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y86     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3380_4 ( .OUT(na3380_2), .IN1(1'b1), .IN2(na633_1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x121y85     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3381_1 ( .OUT(na3381_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(na1962_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x138y93     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3383_1 ( .OUT(na3383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na794_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3383_4 ( .OUT(na3383_2), .IN1(na26_2), .IN2(1'b1), .IN3(na698_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x136y81     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3385_4 ( .OUT(na3385_2), .IN1(na1963_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y85     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3386_4 ( .OUT(na3386_2), .IN1(na634_1), .IN2(~na4170_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x137y92     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3388_1 ( .OUT(na3388_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na795_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3388_4 ( .OUT(na3388_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na699_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y78     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3390_4 ( .OUT(na3390_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1964_1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x127y81     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3391_1 ( .OUT(na3391_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na16_2), .IN6(1'b1), .IN7(1'b1), .IN8(na635_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x131y90     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3393_1 ( .OUT(na3393_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na796_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3393_4 ( .OUT(na3393_2), .IN1(na26_2), .IN2(1'b1), .IN3(na700_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x130y80     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3395_4 ( .OUT(na3395_2), .IN1(1'b1), .IN2(na636_1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x117y77     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3396_1 ( .OUT(na3396_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1965_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x123y88     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3398_1 ( .OUT(na3398_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na701_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3398_4 ( .OUT(na3398_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na797_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x118y75     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3400_4 ( .OUT(na3400_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(na637_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y77     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3401_1 ( .OUT(na3401_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(na1966_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x115y68     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3403_1 ( .OUT(na3403_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(na702_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3403_4 ( .OUT(na3403_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na798_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y66     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3405_1 ( .OUT(na3405_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na638_1), .IN8(na4169_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y65     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3406_1 ( .OUT(na3406_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1967_2), .IN6(na4170_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x132y72     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3408_1 ( .OUT(na3408_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na799_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3408_4 ( .OUT(na3408_2), .IN1(na26_2), .IN2(1'b1), .IN3(na703_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x120y67     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3410_4 ( .OUT(na3410_2), .IN1(1'b1), .IN2(1'b1), .IN3(na639_1), .IN4(na4169_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y67     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3411_1 ( .OUT(na3411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1968_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x121y87     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3413_1 ( .OUT(na3413_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na800_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3413_4 ( .OUT(na3413_2), .IN1(na26_2), .IN2(1'b1), .IN3(na704_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y79     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3415_4 ( .OUT(na3415_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(na640_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y81     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3416_1 ( .OUT(na3416_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3237_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x128y90     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3418_1 ( .OUT(na3418_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na801_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3418_4 ( .OUT(na3418_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na705_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y82     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3420_4 ( .OUT(na3420_2), .IN1(1'b1), .IN2(na641_1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x107y77     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3421_4 ( .OUT(na3421_2), .IN1(na16_2), .IN2(na3238_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x127y91     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3423_1 ( .OUT(na3423_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(1'b1), .IN8(na706_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3423_4 ( .OUT(na3423_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na802_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y95     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3425_1 ( .OUT(na3425_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3239_1), .IN7(1'b1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y87     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3426_4 ( .OUT(na3426_2), .IN1(~na16_2), .IN2(1'b1), .IN3(1'b1), .IN4(na642_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x114y84     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3428_1 ( .OUT(na3428_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(1'b1), .IN8(na707_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3428_4 ( .OUT(na3428_2), .IN1(na26_1), .IN2(1'b1), .IN3(na803_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y80     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3430_1 ( .OUT(na3430_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na643_1), .IN6(1'b1), .IN7(na15_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x107y78     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3431_4 ( .OUT(na3431_2), .IN1(na16_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3240_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x111y81     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3433_1 ( .OUT(na3433_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na804_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3433_4 ( .OUT(na3433_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na708_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y79     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3435_1 ( .OUT(na3435_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na15_2), .IN8(na644_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y77     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3436_4 ( .OUT(na3436_2), .IN1(na16_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3241_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y83     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3438_1 ( .OUT(na3438_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na805_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3438_4 ( .OUT(na3438_2), .IN1(na26_2), .IN2(na709_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y78     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3440_1 ( .OUT(na3440_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na15_2), .IN8(na645_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y73     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3441_4 ( .OUT(na3441_2), .IN1(na16_2), .IN2(na3242_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x107y69     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3443_1 ( .OUT(na3443_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(na710_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3443_4 ( .OUT(na3443_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na806_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y66     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3445_1 ( .OUT(na3445_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3243_1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y68     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3446_4 ( .OUT(na3446_2), .IN1(~na16_2), .IN2(1'b1), .IN3(1'b1), .IN4(na646_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x109y69     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3448_1 ( .OUT(na3448_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na807_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3448_4 ( .OUT(na3448_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na711_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x120y65     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3450_4 ( .OUT(na3450_2), .IN1(na3244_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y67     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3451_4 ( .OUT(na3451_2), .IN1(~na16_2), .IN2(na647_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y69     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3453_1 ( .OUT(na3453_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na241_1), .IN7(na240_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x80y95     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3454_4 ( .OUT(na3454_2), .IN1(~na234_1), .IN2(~na1814_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x86y94     80'h00_0078_00_0000_0C66_AC9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3456_1 ( .OUT(na3456_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na223_2), .IN7(na225_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3456_4 ( .OUT(na3456_2), .IN1(na1162_1), .IN2(1'b0), .IN3(na1160_1), .IN4(~na1164_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x87y93     80'h00_0078_00_0000_0C66_9069
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3457_1 ( .OUT(na3457_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1160_1), .IN8(~na1156_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3457_4 ( .OUT(na3457_2), .IN1(na1162_1), .IN2(~na1151_1), .IN3(na1160_1), .IN4(na1164_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y95     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3459_1 ( .OUT(na3459_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na227_1), .IN7(1'b1), .IN8(na4106_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y91     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3460_4 ( .OUT(na3460_2), .IN1(1'b1), .IN2(1'b1), .IN3(na225_1), .IN4(~na3456_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x85y93     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3463_1 ( .OUT(na3463_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1160_1), .IN8(~na1164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y92     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3466_1 ( .OUT(na3466_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1811_1), .IN6(na1814_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y86     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3467_1 ( .OUT(na3467_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na246_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na248_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x80y96     80'h00_0060_00_0000_0C06_FFA5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3468_4 ( .OUT(na3468_2), .IN1(~na234_1), .IN2(1'b0), .IN3(na4360_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y82     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3469_1 ( .OUT(na3469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1811_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na228_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x85y91     80'h00_0078_00_0000_0C66_CA09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3470_1 ( .OUT(na3470_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na244_1), .IN6(1'b0), .IN7(1'b0), .IN8(na3456_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3470_4 ( .OUT(na3470_2), .IN1(~na1162_1), .IN2(na1166_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x83y91     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3471_4 ( .OUT(na3471_2), .IN1(1'b0), .IN2(1'b0), .IN3(na225_2), .IN4(na4106_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y90     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3472_1 ( .OUT(na3472_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na242_2), .IN8(~na253_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x81y88     80'h00_0078_00_0000_0C88_CA1F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3475_1 ( .OUT(na3475_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na244_1), .IN6(1'b1), .IN7(1'b1), .IN8(na4106_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3475_4 ( .OUT(na3475_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na225_2), .IN4(~na245_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x87y90     80'h00_0078_00_0000_0C66_096A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3477_1 ( .OUT(na3477_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na244_1), .IN6(~na1151_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3477_4 ( .OUT(na3477_2), .IN1(na3470_2), .IN2(1'b0), .IN3(na1160_1), .IN4(na1156_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x85y83     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3478_4 ( .OUT(na3478_2), .IN1(1'b0), .IN2(1'b0), .IN3(na240_2), .IN4(~na248_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x129y76     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3480_4 ( .OUT(na3480_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2099_2), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y73     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3481_4 ( .OUT(na3481_2), .IN1(~na16_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2355_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x80y83     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3485_1 ( .OUT(na3485_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na246_1), .IN6(na241_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x81y91     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3487_4 ( .OUT(na3487_2), .IN1(1'b0), .IN2(1'b0), .IN3(na240_2), .IN4(na4380_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x139y79     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3489_1 ( .OUT(na3489_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2100_1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y71     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3490_4 ( .OUT(na3490_2), .IN1(na2356_1), .IN2(~na4170_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x130y69     80'h00_0018_00_0000_0C88_7AFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3494_1 ( .OUT(na3494_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na282_1), .IN6(1'b0), .IN7(~na15_2), .IN8(~na2357_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y85     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3496_1 ( .OUT(na3496_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na16_2), .IN6(1'b1), .IN7(na2101_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x134y72     80'h00_0060_00_0000_0C08_FF3D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3497_4 ( .OUT(na3497_2), .IN1(~na21_1), .IN2(na3500_1), .IN3(1'b0), .IN4(~na284_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y80     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3500_1 ( .OUT(na3500_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2412_2), .IN8(~na1144_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y91     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3501_1 ( .OUT(na3501_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na225_2), .IN8(na253_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x89y88     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3502_1 ( .OUT(na3502_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na242_2), .IN8(~na4106_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y65     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3504_4 ( .OUT(na3504_2), .IN1(1'b1), .IN2(na2102_1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y68     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3505_1 ( .OUT(na3505_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na16_2), .IN6(1'b1), .IN7(na2358_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x129y70     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3509_4 ( .OUT(na3509_2), .IN1(1'b1), .IN2(na2103_2), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y69     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3510_4 ( .OUT(na3510_2), .IN1(~na16_2), .IN2(na2359_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y65     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3515_1 ( .OUT(na3515_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na16_2), .IN6(1'b1), .IN7(na2360_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y63     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3519_4 ( .OUT(na3519_2), .IN1(1'b1), .IN2(na2361_2), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x120y64     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3520_1 ( .OUT(na3520_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2105_2), .IN6(na4170_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x140y61     80'h00_0060_00_0000_0C08_FF7A
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3524_4 ( .OUT(na3524_2), .IN1(na319_1), .IN2(1'b0), .IN3(~na15_2), .IN4(~na2362_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y61     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3526_4 ( .OUT(na3526_2), .IN1(na2106_2), .IN2(na4170_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x125y66     80'h00_0060_00_0000_0C08_FF3D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3527_4 ( .OUT(na3527_2), .IN1(~na21_1), .IN2(na3530_1), .IN3(1'b0), .IN4(~na321_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y66     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3530_1 ( .OUT(na3530_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1149_2), .IN8(~na2417_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x129y79     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3531_1 ( .OUT(na3531_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1053_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3531_4 ( .OUT(na3531_2), .IN1(na26_2), .IN2(na816_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x124y84     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3536_1 ( .OUT(na3536_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(na862_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3536_4 ( .OUT(na3536_2), .IN1(na1054_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4177_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x139y80     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3541_1 ( .OUT(na3541_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na876_1), .IN7(na349_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x127y79     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3543_4 ( .OUT(na3543_2), .IN1(~na26_2), .IN2(~na871_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x140y81     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3544_1 ( .OUT(na3544_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2404_2), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3544_4 ( .OUT(na3544_2), .IN1(na1055_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4177_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x137y70     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3548_4 ( .OUT(na3548_2), .IN1(1'b1), .IN2(1'b1), .IN3(na349_2), .IN4(na2405_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x137y71     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3550_4 ( .OUT(na3550_2), .IN1(~na26_1), .IN2(~na1056_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x140y74     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3551_1 ( .OUT(na3551_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na349_1), .IN8(na882_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3551_4 ( .OUT(na3551_2), .IN1(na26_2), .IN2(na877_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x125y77     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3555_1 ( .OUT(na3555_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(1'b1), .IN8(na883_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3555_4 ( .OUT(na3555_2), .IN1(na26_1), .IN2(na1057_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x137y67     80'h00_0018_00_0000_0888_5132
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3560_1 ( .OUT(na3560_1), .IN1(na3562_2), .IN2(~na3563_2), .IN3(1'b1), .IN4(~na3561_1), .IN5(~na379_1), .IN6(~na3563_1), .IN7(~na378_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x126y74     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3561_1 ( .OUT(na3561_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(na887_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x131y69     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3562_4 ( .OUT(na3562_2), .IN1(~na26_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1058_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x141y72     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3563_1 ( .OUT(na3563_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2407_1), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3563_4 ( .OUT(na3563_2), .IN1(1'b1), .IN2(1'b1), .IN3(na349_1), .IN4(na889_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x138y69     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3569_1 ( .OUT(na3569_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2408_2), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x136y72     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3571_4 ( .OUT(na3571_2), .IN1(~na26_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1059_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x137y69     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3572_1 ( .OUT(na3572_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na891_1), .IN7(na349_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3572_4 ( .OUT(na3572_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na890_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x117y65     80'h00_0018_00_0000_0888_7BDD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3576_1 ( .OUT(na3576_1), .IN1(~na2114_1), .IN2(na4175_2), .IN3(~na2018_1), .IN4(na25_2), .IN5(na21_2), .IN6(~na1986_1), .IN7(~na2050_1),
                      .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x134y68     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3577_1 ( .OUT(na3577_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na892_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x133y69     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3579_1 ( .OUT(na3579_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na26_1), .IN6(~na1060_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x139y70     80'h00_0078_00_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3580_1 ( .OUT(na3580_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na349_1), .IN8(na894_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3580_4 ( .OUT(na3580_2), .IN1(na2409_1), .IN2(1'b1), .IN3(na349_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y79     80'h00_0018_00_0000_0888_7BDD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3585_1 ( .OUT(na3585_1), .IN1(~na2067_2), .IN2(na4175_2), .IN3(~na2003_2), .IN4(na25_2), .IN5(na21_2), .IN6(~na1971_2), .IN7(~na2035_2),
                      .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y86     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3586_1 ( .OUT(na3586_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na349_1), .IN8(na939_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x145y96     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3588_4 ( .OUT(na3588_2), .IN1(~na2934_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na4178_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x151y93     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3589_1 ( .OUT(na3589_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na349_2), .IN8(na895_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3589_4 ( .OUT(na3589_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1061_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x144y92     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3594_1 ( .OUT(na3594_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(na1062_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3594_4 ( .OUT(na3594_2), .IN1(na26_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2935_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x149y93     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3599_1 ( .OUT(na3599_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na349_2), .IN8(na949_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x149y92     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3601_4 ( .OUT(na3601_2), .IN1(~na26_2), .IN2(1'b0), .IN3(~na2936_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x150y85     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3602_1 ( .OUT(na3602_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na954_1), .IN7(na349_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3602_4 ( .OUT(na3602_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1063_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x153y92     80'h00_0018_00_0000_0888_131C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3606_1 ( .OUT(na3606_1), .IN1(1'b1), .IN2(na3608_2), .IN3(~na3607_1), .IN4(~na3609_2), .IN5(1'b1), .IN6(~na430_1), .IN7(~na431_1),
                      .IN8(~na3609_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y87     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3607_1 ( .OUT(na3607_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na2937_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x141y90     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3608_4 ( .OUT(na3608_2), .IN1(~na26_1), .IN2(1'b0), .IN3(~na1064_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x150y86     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3609_1 ( .OUT(na3609_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na955_2), .IN6(1'b1), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3609_4 ( .OUT(na3609_2), .IN1(na961_1), .IN2(1'b1), .IN3(na349_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x149y83     80'h00_0018_00_0000_0888_321F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3614_1 ( .OUT(na3614_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na439_1), .IN4(~na3619_1), .IN5(na437_1), .IN6(~na440_1), .IN7(1'b1),
                      .IN8(~na3619_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x146y84     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3619_1 ( .OUT(na3619_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(1'b1), .IN7(na2938_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3619_4 ( .OUT(na3619_2), .IN1(na1065_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4177_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x110y71     80'h00_0018_00_0000_0888_7BDD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3621_1 ( .OUT(na3621_1), .IN1(~na2072_1), .IN2(na4175_2), .IN3(~na2008_1), .IN4(na25_2), .IN5(na21_2), .IN6(~na1976_1), .IN7(~na2040_1),
                      .IN8(~na4172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x150y87     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3622_4 ( .OUT(na3622_2), .IN1(1'b1), .IN2(na967_1), .IN3(na349_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x149y84     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3624_1 ( .OUT(na3624_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na26_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na2939_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x151y83     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3625_1 ( .OUT(na3625_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na965_2), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3625_4 ( .OUT(na3625_2), .IN1(na26_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1066_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y86     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3630_4 ( .OUT(na3630_2), .IN1(1'b1), .IN2(na968_2), .IN3(na349_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x146y81     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3632_1 ( .OUT(na3632_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na26_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na2940_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x143y80     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3633_1 ( .OUT(na3633_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na969_1), .IN7(na349_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3633_4 ( .OUT(na3633_2), .IN1(na1067_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4177_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y73     80'h00_0018_00_0000_0888_114F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3637_1 ( .OUT(na3637_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na3640_2), .IN4(na3639_1), .IN5(~na465_1), .IN6(~na3638_2), .IN7(~na3640_1),
                      .IN8(~na466_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y80     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3638_4 ( .OUT(na3638_2), .IN1(na26_2), .IN2(1'b1), .IN3(na2941_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x142y78     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3639_1 ( .OUT(na3639_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na26_1), .IN6(1'b0), .IN7(~na1068_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x146y73     80'h00_0078_00_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3640_1 ( .OUT(na3640_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na970_2), .IN6(1'b1), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3640_4 ( .OUT(na3640_2), .IN1(1'b1), .IN2(na971_1), .IN3(na349_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x142y88     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3646_1 ( .OUT(na3646_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_2), .IN6(na2363_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3646_4 ( .OUT(na3646_2), .IN1(na26_1), .IN2(1'b1), .IN3(na1069_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y82     80'h00_0018_00_0000_0888_315C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3651_1 ( .OUT(na3651_1), .IN1(1'b1), .IN2(na481_2), .IN3(~na4383_2), .IN4(1'b1), .IN5(~na484_1), .IN6(~na3656_2), .IN7(1'b1),
                      .IN8(~na483_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x147y84     80'h00_0078_00_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3656_1 ( .OUT(na3656_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1029_1), .IN7(na349_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3656_4 ( .OUT(na3656_2), .IN1(na2927_1), .IN2(1'b1), .IN3(na349_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x135y86     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3657_1 ( .OUT(na3657_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1070_1), .IN8(~na2364_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x145y91     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3659_4 ( .OUT(na3659_2), .IN1(1'b1), .IN2(1'b1), .IN3(na349_2), .IN4(na2928_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x141y89     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3661_1 ( .OUT(na3661_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2365_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na4178_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x148y82     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3662_1 ( .OUT(na3662_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na349_1), .IN8(na1034_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3662_4 ( .OUT(na3662_2), .IN1(na26_1), .IN2(na1071_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x144y87     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3666_4 ( .OUT(na3666_2), .IN1(na2929_1), .IN2(1'b1), .IN3(na349_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x139y83     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3668_4 ( .OUT(na3668_2), .IN1(~na26_1), .IN2(1'b0), .IN3(~na1072_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x141y82     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3669_1 ( .OUT(na3669_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4196_2), .IN6(1'b1), .IN7(na1040_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3669_4 ( .OUT(na3669_2), .IN1(na26_2), .IN2(na2366_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x147y82     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3673_1 ( .OUT(na3673_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1044_1), .IN7(na349_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3673_4 ( .OUT(na3673_2), .IN1(1'b1), .IN2(1'b1), .IN3(na349_2), .IN4(na2930_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y85     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3675_1 ( .OUT(na3675_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1073_1), .IN6(~na2367_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y80     80'h00_0018_00_0000_0888_112F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3679_1 ( .OUT(na3679_1), .IN1(1'b1), .IN2(1'b1), .IN3(na3681_1), .IN4(~na3682_2), .IN5(~na519_1), .IN6(~na520_1), .IN7(~na3680_2),
                      .IN8(~na3682_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x132y83     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3680_4 ( .OUT(na3680_2), .IN1(na2368_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4178_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x136y81     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3681_1 ( .OUT(na3681_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na26_1), .IN6(1'b0), .IN7(~na1074_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x142y82     80'h00_0078_00_0000_0C88_8F8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3682_1 ( .OUT(na3682_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na349_1), .IN8(na1048_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3682_4 ( .OUT(na3682_2), .IN1(1'b1), .IN2(1'b1), .IN3(na349_2), .IN4(na2931_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x138y70     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3688_4 ( .OUT(na3688_2), .IN1(na26_2), .IN2(1'b1), .IN3(na2369_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x140y77     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3690_1 ( .OUT(na3690_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na26_1), .IN6(1'b0), .IN7(~na1075_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x141y74     80'h00_0078_00_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3691_1 ( .OUT(na3691_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2932_2), .IN6(1'b1), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3691_4 ( .OUT(na3691_2), .IN1(1'b1), .IN2(1'b1), .IN3(na349_1), .IN4(na1050_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x138y76     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3695_1 ( .OUT(na3695_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na26_1), .IN6(1'b1), .IN7(na1076_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3695_4 ( .OUT(na3695_2), .IN1(na26_2), .IN2(na2370_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y66     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3700_4 ( .OUT(na3700_2), .IN1(~na1331_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y59     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3701_1 ( .OUT(na3701_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na548_2), .IN6(1'b1), .IN7(1'b1), .IN8(na547_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x141y59     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3702_1 ( .OUT(na3702_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na539_1), .IN6(~na541_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x82y99     80'h00_0078_00_0000_0C66_CA9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3705_1 ( .OUT(na3705_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3723_2), .IN6(1'b0), .IN7(1'b0), .IN8(na839_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3705_4 ( .OUT(na3705_2), .IN1(na825_1), .IN2(1'b0), .IN3(~na842_2), .IN4(na4247_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y95     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3706_1 ( .OUT(na3706_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1844_1), .IN8(na836_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x91y101     80'h00_0078_00_0000_0C66_3AA5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3711_1 ( .OUT(na3711_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na825_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1172_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3711_4 ( .OUT(na3711_2), .IN1(~na1178_1), .IN2(1'b0), .IN3(na1182_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y100     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3715_1 ( .OUT(na3715_1), .IN1(1'b1), .IN2(na827_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4322_2), .IN8(~na1172_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x89y100     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3716_4 ( .OUT(na3716_2), .IN1(na825_1), .IN2(1'b0), .IN3(na824_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x80y96     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3717_1 ( .OUT(na3717_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1842_1), .IN6(1'b0), .IN7(na1844_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x85y97     80'h00_0060_00_0000_0C06_FF5C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3718_4 ( .OUT(na3718_2), .IN1(1'b0), .IN2(na846_2), .IN3(~na848_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x80y101     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3719_1 ( .OUT(na3719_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na829_1), .IN7(1'b0), .IN8(na836_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x79y102     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3720_4 ( .OUT(na3720_2), .IN1(~na1842_1), .IN2(1'b0), .IN3(1'b0), .IN4(na836_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y99     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3721_1 ( .OUT(na3721_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na822_2), .IN7(1'b0), .IN8(na4257_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x85y98     80'h00_0060_00_0000_0C06_FFC3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3722_4 ( .OUT(na3722_2), .IN1(1'b0), .IN2(~na827_1), .IN3(1'b0), .IN4(na839_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x81y97     80'h00_0078_00_0000_0C66_C309
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3723_1 ( .OUT(na3723_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na820_1), .IN7(1'b0), .IN8(na839_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3723_4 ( .OUT(na3723_2), .IN1(~na825_1), .IN2(na827_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y95     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3724_1 ( .OUT(na3724_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na854_1), .IN6(1'b0), .IN7(na842_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x88y102     80'h00_0078_00_0000_0C66_0990
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3728_1 ( .OUT(na3728_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1168_1), .IN6(na844_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3728_4 ( .OUT(na3728_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na824_1), .IN4(na4386_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x84y100     80'h00_0060_00_0000_0C06_FFA5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3729_4 ( .OUT(na3729_2), .IN1(~na3723_2), .IN2(1'b0), .IN3(na848_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y80     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3730_1 ( .OUT(na3730_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3256_1), .IN7(na70_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x89y98     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3732_4 ( .OUT(na3732_2), .IN1(na3723_2), .IN2(1'b0), .IN3(1'b0), .IN4(na3728_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y94     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3734_1 ( .OUT(na3734_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na846_2), .IN7(na3705_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y84     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3735_1 ( .OUT(na3735_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na76_1), .IN7(na3257_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y83     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3736_1 ( .OUT(na3736_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3258_1), .IN6(1'b0), .IN7(1'b0), .IN8(na82_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x88y96     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3737_4 ( .OUT(na3737_2), .IN1(na854_1), .IN2(~na827_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x92y98     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3738_1 ( .OUT(na3738_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na827_1), .IN7(na842_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y71     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3739_4 ( .OUT(na3739_2), .IN1(1'b0), .IN2(na3259_1), .IN3(na88_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y77     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3740_1 ( .OUT(na3740_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na94_1), .IN6(1'b0), .IN7(1'b0), .IN8(na3260_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x117y75     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3741_4 ( .OUT(na3741_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3261_1), .IN4(na100_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x119y70     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3742_4 ( .OUT(na3742_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3262_1), .IN4(na106_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x118y68     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3743_4 ( .OUT(na3743_2), .IN1(na3263_1), .IN2(1'b0), .IN3(1'b0), .IN4(na112_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x149y99     80'h00_0078_00_0000_0C66_90A3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3744_1 ( .OUT(na3744_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1184_1), .IN8(na917_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3744_4 ( .OUT(na3744_2), .IN1(1'b0), .IN2(~na900_1), .IN3(na3766_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x151y102     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3745_1 ( .OUT(na3745_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3759_2), .IN8(na911_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x144y104     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3750_4 ( .OUT(na3750_2), .IN1(1'b0), .IN2(na900_1), .IN3(1'b0), .IN4(na899_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x147y101     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3752_1 ( .OUT(na3752_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na901_1), .IN8(na899_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x137y101     80'h00_0078_00_0000_0C66_5CC9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3753_1 ( .OUT(na3753_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na900_1), .IN7(~na1184_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3753_4 ( .OUT(na3753_2), .IN1(na1192_1), .IN2(~na1196_1), .IN3(1'b0), .IN4(na1194_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x154y102     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3756_4 ( .OUT(na3756_2), .IN1(na906_1), .IN2(1'b0), .IN3(na3759_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x154y100     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3757_1 ( .OUT(na3757_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4405_2), .IN6(na929_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x153y101     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3758_1 ( .OUT(na3758_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1847_2), .IN7(na3759_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x148y101     80'h00_0078_00_0000_0C66_CCC6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3759_1 ( .OUT(na3759_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1847_2), .IN7(1'b0), .IN8(na911_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3759_4 ( .OUT(na3759_2), .IN1(na1848_1), .IN2(na915_2), .IN3(1'b0), .IN4(na916_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x149y98     80'h00_0078_00_0000_0C88_CCF4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3763_1 ( .OUT(na3763_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na929_2), .IN7(1'b1), .IN8(na917_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3763_4 ( .OUT(na3763_2), .IN1(~na920_1), .IN2(na929_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x149y103     80'h00_0078_00_0000_0C66_A3C9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3765_1 ( .OUT(na3765_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3768_2), .IN7(na921_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3765_4 ( .OUT(na3765_2), .IN1(~na932_1), .IN2(na900_1), .IN3(1'b0), .IN4(na899_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x140y101     80'h00_0078_00_0000_0C66_CA90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3766_1 ( .OUT(na3766_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3753_2), .IN6(1'b0), .IN7(1'b0), .IN8(na917_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3766_4 ( .OUT(na3766_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1198_1), .IN4(~na1194_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x149y97     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3767_1 ( .OUT(na3767_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na901_1), .IN8(na4277_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x149y100     80'h00_0078_00_0000_0C66_9090
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3768_1 ( .OUT(na3768_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na921_1), .IN8(~na898_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3768_4 ( .OUT(na3768_2), .IN1(1'b0), .IN2(1'b0), .IN3(na901_1), .IN4(~na899_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x146y97     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3769_4 ( .OUT(na3769_2), .IN1(na932_1), .IN2(~na938_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x149y96     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3770_1 ( .OUT(na3770_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na118_1), .IN7(1'b0), .IN8(na3264_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x155y99     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3771_4 ( .OUT(na3771_2), .IN1(1'b0), .IN2(na929_1), .IN3(na4280_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x151y99     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3772_1 ( .OUT(na3772_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3744_2), .IN6(na3768_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x153y97     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3774_4 ( .OUT(na3774_2), .IN1(na3765_2), .IN2(na929_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y96     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3775_1 ( .OUT(na3775_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3265_1), .IN8(na124_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x155y92     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3776_4 ( .OUT(na3776_2), .IN1(na130_1), .IN2(1'b0), .IN3(na3266_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x144y100     80'h00_0018_00_0000_0C66_5C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3777_1 ( .OUT(na3777_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na938_1), .IN7(~na901_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x149y101     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3778_4 ( .OUT(na3778_2), .IN1(na932_1), .IN2(1'b0), .IN3(~na901_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x147y90     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3779_1 ( .OUT(na3779_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3267_1), .IN8(na136_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x143y93     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3780_4 ( .OUT(na3780_2), .IN1(na3268_1), .IN2(1'b0), .IN3(na142_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x140y92     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3781_4 ( .OUT(na3781_2), .IN1(1'b0), .IN2(na3269_1), .IN3(na148_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x142y78     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3782_4 ( .OUT(na3782_2), .IN1(na3270_1), .IN2(1'b0), .IN3(1'b0), .IN4(na154_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x146y77     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3783_1 ( .OUT(na3783_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na160_1), .IN6(1'b0), .IN7(1'b0), .IN8(na3271_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x92y103     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3786_4 ( .OUT(na3786_2), .IN1(1'b0), .IN2(na984_1), .IN3(1'b0), .IN4(na3800_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x97y99     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3790_1 ( .OUT(na3790_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na979_1), .IN7(1'b0), .IN8(na978_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x103y102     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3792_4 ( .OUT(na3792_2), .IN1(na977_1), .IN2(1'b1), .IN3(1'b1), .IN4(na978_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x104y98     80'h00_0078_00_0000_0C66_099A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3793_1 ( .OUT(na3793_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1200_1), .IN6(na979_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3793_4 ( .OUT(na3793_2), .IN1(na1210_1), .IN2(1'b0), .IN3(~na1212_1), .IN4(na1208_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x91y102     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3796_1 ( .OUT(na3796_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1852_1), .IN6(1'b0), .IN7(1'b0), .IN8(na3800_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x93y101     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3798_1 ( .OUT(na3798_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na989_1), .IN8(na3800_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x96y100     80'h00_0078_00_0000_0C66_5AA6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3800_1 ( .OUT(na3800_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1852_1), .IN6(1'b0), .IN7(~na989_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3800_4 ( .OUT(na3800_2), .IN1(na1853_1), .IN2(na994_1), .IN3(na993_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x99y101     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3801_1 ( .OUT(na3801_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1002_2), .IN6(na1001_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x104y100     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3802_4 ( .OUT(na3802_2), .IN1(~na1007_1), .IN2(na1005_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x103y100     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3804_1 ( .OUT(na3804_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na977_2), .IN6(1'b0), .IN7(1'b0), .IN8(na4288_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x109y103     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3806_4 ( .OUT(na3806_2), .IN1(na1003_1), .IN2(1'b0), .IN3(~na1013_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x102y102     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3808_1 ( .OUT(na3808_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1007_1), .IN6(~na1001_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y83     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3809_4 ( .OUT(na3809_2), .IN1(1'b0), .IN2(na3272_1), .IN3(1'b0), .IN4(na166_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x100y98     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3811_4 ( .OUT(na3811_2), .IN1(1'b0), .IN2(na1001_2), .IN3(na1006_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x108y102     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3813_4 ( .OUT(na3813_2), .IN1(na1002_2), .IN2(na1005_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x135y89     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3814_1 ( .OUT(na3814_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3273_1), .IN8(na172_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x133y90     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3815_4 ( .OUT(na3815_2), .IN1(na3274_1), .IN2(na178_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x100y99     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3816_1 ( .OUT(na3816_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na977_2), .IN6(1'b0), .IN7(na1013_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x109y92     80'h00_0060_00_0000_0C06_FF3A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3817_4 ( .OUT(na3817_2), .IN1(na1003_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na4288_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x134y87     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3818_1 ( .OUT(na3818_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3275_1), .IN7(na184_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y86     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3819_1 ( .OUT(na3819_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na190_1), .IN7(1'b0), .IN8(na3276_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y84     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3820_1 ( .OUT(na3820_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3277_1), .IN6(1'b0), .IN7(na196_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x129y78     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3821_1 ( .OUT(na3821_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na202_1), .IN6(1'b0), .IN7(na3278_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x128y74     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3822_4 ( .OUT(na3822_2), .IN1(1'b0), .IN2(na208_1), .IN3(na3279_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x105y95     80'h00_0078_00_0000_0C66_6006
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3871_1 ( .OUT(na3871_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3248_1), .IN8(na13_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3871_4 ( .OUT(na3871_2), .IN1(na3294_2), .IN2(na1859_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x128y77     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3872_1 ( .OUT(na3872_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na27_1), .IN8(na3249_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y78     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3873_4 ( .OUT(na3873_2), .IN1(na34_1), .IN2(1'b0), .IN3(1'b0), .IN4(na3250_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x125y67     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3874_1 ( .OUT(na3874_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na40_1), .IN6(na3251_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x117y69     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3875_4 ( .OUT(na3875_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3252_1), .IN4(na46_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y69     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3876_4 ( .OUT(na3876_2), .IN1(na3253_1), .IN2(1'b0), .IN3(1'b0), .IN4(na52_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y66     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3877_1 ( .OUT(na3877_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na58_1), .IN6(1'b0), .IN7(1'b0), .IN8(na3254_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x116y67     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3878_4 ( .OUT(na3878_2), .IN1(1'b0), .IN2(na64_1), .IN3(1'b0), .IN4(na3255_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x153y81     80'h00_0018_00_0000_0888_2A1C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3952_1 ( .OUT(na3952_1), .IN1(1'b1), .IN2(na3955_2), .IN3(~na3954_1), .IN4(~na3956_2), .IN5(na3953_2), .IN6(1'b1), .IN7(na1233_1),
                      .IN8(~na1230_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x155y89     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3953_4 ( .OUT(na3953_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1117_1), .IN4(~na1222_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x152y81     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3954_1 ( .OUT(na3954_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1017_1), .IN8(na1224_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x149y80     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3955_4 ( .OUT(na3955_2), .IN1(~na1245_2), .IN2(1'b0), .IN3(~na1141_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x146y82     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3956_4 ( .OUT(na3956_2), .IN1(1'b1), .IN2(na1229_1), .IN3(1'b1), .IN4(na1101_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x153y75     80'h00_0018_00_0000_0888_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3958_1 ( .OUT(na3958_1), .IN1(~na1319_1), .IN2(~na1286_1), .IN3(~na1297_1), .IN4(~na1857_1), .IN5(~na1253_1), .IN6(~na1265_1),
                      .IN7(~na1308_1), .IN8(~na1219_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x152y84     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3959_1 ( .OUT(na3959_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1069_1), .IN8(~na1235_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x151y86     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3960_4 ( .OUT(na3960_2), .IN1(na1093_1), .IN2(na4332_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x149y80     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3961_1 ( .OUT(na3961_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1238_2), .IN8(~na1053_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x153y91     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3962_4 ( .OUT(na3962_2), .IN1(1'b1), .IN2(na1251_2), .IN3(na1085_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x155y87     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3963_1 ( .OUT(na3963_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1243_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na939_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x152y80     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3964_4 ( .OUT(na3964_2), .IN1(na1243_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2918_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x148y75     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3965_1 ( .OUT(na3965_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1245_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1133_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x148y77     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3966_1 ( .OUT(na3966_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1077_1), .IN7(na1246_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x154y88     80'h00_0078_00_0000_0CEE_5533
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3967_1 ( .OUT(na3967_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1236_2), .IN6(1'b0), .IN7(~na1125_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3967_4 ( .OUT(na3967_2), .IN1(1'b0), .IN2(~na1251_1), .IN3(1'b0), .IN4(~na1061_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y77     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3968_1 ( .OUT(na3968_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1109_1), .IN8(na1224_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x149y78     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3970_1 ( .OUT(na3970_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na861_1), .IN8(na1235_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y84     80'h00_0018_00_0000_0888_8841
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3971_1 ( .OUT(na3971_1), .IN1(~na3973_2), .IN2(~na3977_2), .IN3(~na3975_2), .IN4(na1259_1), .IN5(na3972_1), .IN6(na3974_2),
                      .IN7(na1258_2), .IN8(na3976_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x153y91     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3972_1 ( .OUT(na3972_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1118_1), .IN7(1'b0), .IN8(~na1222_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y79     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3973_4 ( .OUT(na3973_2), .IN1(1'b1), .IN2(na1229_1), .IN3(1'b1), .IN4(na1102_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x149y84     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3974_4 ( .OUT(na3974_2), .IN1(~na1054_1), .IN2(1'b0), .IN3(~na1238_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x152y79     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3975_4 ( .OUT(na3975_2), .IN1(na1243_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2919_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x152y82     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3976_1 ( .OUT(na3976_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1029_1), .IN7(1'b0), .IN8(~na1224_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x151y88     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3977_4 ( .OUT(na3977_2), .IN1(na1236_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1094_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x154y91     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3983_1 ( .OUT(na3983_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1086_1), .IN6(na1251_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x154y87     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3984_4 ( .OUT(na3984_2), .IN1(~na1126_1), .IN2(~na4333_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x153y90     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3985_1 ( .OUT(na3985_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1243_2), .IN6(na948_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x151y78     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3986_1 ( .OUT(na3986_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1229_1), .IN7(~na1103_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x151y87     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3987_4 ( .OUT(na3987_2), .IN1(na1236_1), .IN2(1'b1), .IN3(na1095_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x152y87     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3988_1 ( .OUT(na3988_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1071_1), .IN7(1'b0), .IN8(~na1235_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x151y80     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3989_4 ( .OUT(na3989_2), .IN1(na1079_1), .IN2(1'b1), .IN3(na1246_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x154y90     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3990_1 ( .OUT(na3990_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1119_1), .IN8(~na1222_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x156y88     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3991_4 ( .OUT(na3991_2), .IN1(1'b1), .IN2(na1251_1), .IN3(1'b1), .IN4(na1063_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x149y79     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3994_1 ( .OUT(na3994_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1055_1), .IN6(1'b0), .IN7(~na1238_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x156y88     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3995_1 ( .OUT(na3995_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1251_2), .IN7(1'b1), .IN8(na1087_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x149y82     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3996_4 ( .OUT(na3996_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1111_1), .IN4(~na1224_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x152y79     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3997_1 ( .OUT(na3997_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2920_2), .IN6(1'b1), .IN7(1'b1), .IN8(na4335_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x152y81     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3998_4 ( .OUT(na3998_2), .IN1(1'b0), .IN2(~na876_1), .IN3(1'b0), .IN4(~na1235_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x153y83     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3999_4 ( .OUT(na3999_2), .IN1(na1243_2), .IN2(na954_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x154y76     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4000_4 ( .OUT(na4000_2), .IN1(~na1245_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na1144_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x153y72     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4001_4 ( .OUT(na4001_2), .IN1(na1245_1), .IN2(na1135_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x149y77     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4003_4 ( .OUT(na4003_2), .IN1(1'b0), .IN2(~na1056_1), .IN3(~na1238_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x150y75     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4005_4 ( .OUT(na4005_2), .IN1(~na1245_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na1145_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x152y86     80'h00_0078_00_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4006_1 ( .OUT(na4006_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1251_2), .IN7(1'b1), .IN8(na1088_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4006_4 ( .OUT(na4006_2), .IN1(1'b1), .IN2(na1251_1), .IN3(na1064_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x151y79     80'h00_0018_00_0000_0888_8812
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4013_1 ( .OUT(na4013_1), .IN1(na1291_1), .IN2(~na1289_1), .IN3(~na4014_1), .IN4(~na4016_2), .IN5(na1291_2), .IN6(na1294_1),
                      .IN7(na1293_2), .IN8(na4015_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y81     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4014_1 ( .OUT(na4014_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1236_1), .IN6(na1097_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x146y74     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4015_1 ( .OUT(na4015_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1057_1), .IN7(~na1238_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x152y84     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4016_4 ( .OUT(na4016_2), .IN1(na1243_2), .IN2(1'b1), .IN3(1'b1), .IN4(na964_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x154y73     80'h00_0078_00_0000_0CEE_3335
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4025_1 ( .OUT(na4025_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1044_1), .IN7(1'b0), .IN8(~na1224_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4025_4 ( .OUT(na4025_2), .IN1(~na1243_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na2922_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x153y70     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4026_1 ( .OUT(na4026_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1245_2), .IN6(1'b1), .IN7(na1146_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x150y74     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4028_4 ( .OUT(na4028_2), .IN1(na1245_1), .IN2(na1137_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x152y77     80'h00_0018_00_0000_0888_8812
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4029_1 ( .OUT(na4029_1), .IN1(na1303_1), .IN2(~na4031_1), .IN3(~na4035_2), .IN4(~na4033_1), .IN5(na4030_1), .IN6(na1302_2),
                      .IN7(na4032_2), .IN8(na4034_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x151y85     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4030_1 ( .OUT(na4030_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1122_1), .IN7(1'b0), .IN8(~na1222_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x153y84     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4031_1 ( .OUT(na4031_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1251_1), .IN7(1'b1), .IN8(na1066_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x148y75     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4032_4 ( .OUT(na4032_2), .IN1(1'b0), .IN2(~na1229_1), .IN3(~na1106_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y80     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4033_1 ( .OUT(na4033_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1236_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x148y78     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4034_4 ( .OUT(na4034_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1114_1), .IN4(~na1224_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x150y77     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4035_4 ( .OUT(na4035_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1238_2), .IN4(na1058_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x151y71     80'h00_0078_00_0000_0CEE_0753
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4041_1 ( .OUT(na4041_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1245_2), .IN6(~na1147_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4041_4 ( .OUT(na4041_2), .IN1(1'b0), .IN2(~na1251_2), .IN3(~na1090_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y69     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4042_4 ( .OUT(na4042_2), .IN1(na1245_1), .IN2(na1138_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y74     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4044_4 ( .OUT(na4044_2), .IN1(1'b1), .IN2(na4337_2), .IN3(na1082_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x149y71     80'h00_0018_00_0000_0888_8841
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4045_1 ( .OUT(na4045_1), .IN1(~na1310_1), .IN2(~na4048_2), .IN3(~na4046_2), .IN4(na1313_1), .IN5(na4047_1), .IN6(na1316_2),
                      .IN7(na1315_1), .IN8(na1313_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x148y77     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4046_4 ( .OUT(na4046_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1075_1), .IN4(na1235_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x153y79     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4047_1 ( .OUT(na4047_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1123_1), .IN7(1'b0), .IN8(~na1222_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x147y76     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4048_4 ( .OUT(na4048_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1115_1), .IN4(na1224_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x150y70     80'h00_0078_00_0000_0CEE_5507
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4057_1 ( .OUT(na4057_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1236_2), .IN6(1'b0), .IN7(~na1131_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4057_4 ( .OUT(na4057_2), .IN1(~na1245_2), .IN2(~na1148_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x151y77     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4058_4 ( .OUT(na4058_2), .IN1(na1236_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1099_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x149y68     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4060_1 ( .OUT(na4060_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1245_1), .IN6(1'b1), .IN7(na1139_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x151y68     80'h00_0018_00_0000_0888_4444
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4061_1 ( .OUT(na4061_1), .IN1(~na4066_1), .IN2(na1326_1), .IN3(~na1323_1), .IN4(na1325_1), .IN5(~na4066_2), .IN6(na4065_1),
                      .IN7(~na1323_2), .IN8(na4063_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x148y76     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4063_4 ( .OUT(na4063_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1076_1), .IN4(~na1235_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x153y78     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4065_1 ( .OUT(na4065_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1124_1), .IN7(1'b0), .IN8(~na1222_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x145y69     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4066_1 ( .OUT(na4066_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1084_1), .IN7(na1246_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4066_4 ( .OUT(na4066_2), .IN1(na1245_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1140_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x147y69     80'h00_0078_00_0000_0CEE_0755
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4072_1 ( .OUT(na4072_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1108_1), .IN6(~na1229_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4072_4 ( .OUT(na4072_2), .IN1(~na1245_2), .IN2(1'b0), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x154y72     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4073_4 ( .OUT(na4073_2), .IN1(na1236_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1132_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x150y74     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4075_1 ( .OUT(na4075_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1236_1), .IN6(na1100_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x116y65     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4076_4 ( .OUT(na4076_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1387_2), .IN4(na1332_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y67     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4077_1 ( .OUT(na4077_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1859_1), .IN7(na1387_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y64     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4078_4 ( .OUT(na4078_2), .IN1(1'b1), .IN2(~na1361_1), .IN3(~na3196_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y60     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4081_4 ( .OUT(na4081_2), .IN1(1'b1), .IN2(~na1348_1), .IN3(na3196_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x85y59     80'h00_0060_00_0000_0C0E_FFE3
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a4084_4 ( .OUT(na4084_2), .IN1(1'b0), .IN2(~na1361_1), .IN3(na3196_2), .IN4(na1338_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x127y75     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4088_4 ( .OUT(na4088_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1142_1), .IN4(~na25_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x134y75     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4089_1 ( .OUT(na4089_1), .IN1(~na552_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4171_2), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x130y80     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4091_1 ( .OUT(na4091_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na552_2), .IN6(1'b1), .IN7(na1142_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y67     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4093_1 ( .OUT(na4093_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1142_1), .IN8(~na1332_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y74     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4103_4 ( .OUT(na4103_2), .IN1(~na16_2), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x140y63     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4104_1 ( .OUT(na4104_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3143_1), .IN7(1'b1), .IN8(~na3145_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x139y63     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4105_4 ( .OUT(na4105_2), .IN1(1'b1), .IN2(na3143_1), .IN3(1'b1), .IN4(na3145_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x88y92     80'h00_0078_00_0000_0C66_CA66
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4106_1 ( .OUT(na4106_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3457_2), .IN6(1'b0), .IN7(1'b0), .IN8(na1156_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4106_4 ( .OUT(na4106_2), .IN1(~na1162_1), .IN2(~na1166_1), .IN3(na1158_1), .IN4(na1156_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y96     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4108_1 ( .OUT(na4108_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1151_1), .IN7(na225_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x87y95     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4109_4 ( .OUT(na4109_2), .IN1(na1162_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1164_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y78     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4112_1 ( .OUT(na4112_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1141_2), .IN8(~na2410_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x130y75     80'h00_0018_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4114_1 ( .OUT(na4114_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_1), .IN6(na4112_1), .IN7(1'b0), .IN8(na1816_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x119y77     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4115_1 ( .OUT(na4115_1), .IN1(~na1987_2), .IN2(1'b0), .IN3(~na2019_2), .IN4(na25_2), .IN5(~na21_1), .IN6(~na2051_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x131y70     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4116_4 ( .OUT(na4116_2), .IN1(1'b1), .IN2(1'b1), .IN3(na214_1), .IN4(~na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y74     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4117_1 ( .OUT(na4117_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2411_1), .IN6(~na1143_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x134y71     80'h00_0018_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4119_1 ( .OUT(na4119_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_1), .IN6(na4117_1), .IN7(1'b0), .IN8(na1821_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x125y81     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4120_1 ( .OUT(na4120_1), .IN1(~na1988_1), .IN2(1'b0), .IN3(~na2020_1), .IN4(na25_2), .IN5(~na21_1), .IN6(~na2052_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x136y69     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4121_4 ( .OUT(na4121_2), .IN1(na264_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1451_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x131y72     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4122_1 ( .OUT(na4122_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2413_1), .IN8(~na1145_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x138y75     80'h00_0018_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4124_1 ( .OUT(na4124_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na21_1), .IN6(na4122_1), .IN7(na1826_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x120y72     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4125_1 ( .OUT(na4125_1), .IN1(~na1990_1), .IN2(1'b0), .IN3(~na2022_1), .IN4(na25_2), .IN5(~na21_1), .IN6(~na2054_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x144y59     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4126_1 ( .OUT(na4126_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na287_1), .IN8(~na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x125y70     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4127_1 ( .OUT(na4127_1), .IN1(1'b1), .IN2(~na1333_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1146_2), .IN8(~na2414_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x128y65     80'h00_0060_00_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4129_4 ( .OUT(na4129_2), .IN1(~na21_1), .IN2(na4127_1), .IN3(na1831_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x117y73     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4130_1 ( .OUT(na4130_1), .IN1(~na1991_2), .IN2(1'b0), .IN3(~na2023_2), .IN4(na25_2), .IN5(~na21_1), .IN6(~na2055_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x127y66     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4131_1 ( .OUT(na4131_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na295_1), .IN8(~na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x139y68     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4133_1 ( .OUT(na4133_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2104_1), .IN8(na1451_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x108y73     80'h00_0018_00_0000_0888_F7D5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a4134_1 ( .OUT(na4134_1), .IN1(~na1992_1), .IN2(1'b0), .IN3(~na2024_1), .IN4(na25_2), .IN5(~na21_1), .IN6(~na2056_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x86y103     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4138_1 ( .OUT(na4138_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4250_2), .IN5(~na825_1), .IN6(1'b0), .IN7(~na824_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y101     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4142_4 ( .OUT(na4142_2), .IN1(na825_1), .IN2(na827_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y102     80'h00_0078_00_0000_0C88_F4C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4143_1 ( .OUT(na4143_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1168_1), .IN6(na822_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4143_4 ( .OUT(na4143_2), .IN1(~na3711_2), .IN2(1'b1), .IN3(1'b1), .IN4(na821_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y102     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4148_1 ( .OUT(na4148_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4288_2), .IN5(1'b0), .IN6(~na979_1), .IN7(1'b0), .IN8(~na978_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x122y70     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4154_1 ( .OUT(na4154_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1859_1), .IN7(1'b1), .IN8(na1858_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x120y69     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4155_1 ( .OUT(na4155_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1859_1), .IN7(1'b1), .IN8(~na1858_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y64     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4156_1 ( .OUT(na4156_1), .IN1(1'b1), .IN2(na1333_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2416_2), .IN6(~na1148_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x129y68     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4157_4 ( .OUT(na4157_2), .IN1(~na21_1), .IN2(na4156_1), .IN3(~na311_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x160y73     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4158_4 ( .OUT(na4158_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1362_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4158_6 ( .RAM_O2(na4158_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4158_2), .COMP_OUT(1'b0) );
// C_///AND/      x107y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4159_4 ( .OUT(na4159_2), .IN1(na3_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4159_6 ( .RAM_O2(na4159_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4159_2), .COMP_OUT(1'b0) );
// C_///AND/      x111y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4160_4 ( .OUT(na4160_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4160_6 ( .RAM_O2(na4160_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4160_2), .COMP_OUT(1'b0) );
// C_///AND/      x115y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4161_4 ( .OUT(na4161_2), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4161_6 ( .RAM_O2(na4161_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4161_2), .COMP_OUT(1'b0) );
// C_///AND/      x119y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4162_4 ( .OUT(na4162_2), .IN1(1'b1), .IN2(na5_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4162_6 ( .RAM_O2(na4162_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4162_2), .COMP_OUT(1'b0) );
// C_///AND/      x123y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4163_4 ( .OUT(na4163_2), .IN1(1'b1), .IN2(na5_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4163_6 ( .RAM_O2(na4163_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4163_2), .COMP_OUT(1'b0) );
// C_///AND/      x127y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4164_4 ( .OUT(na4164_2), .IN1(na6_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4164_6 ( .RAM_O2(na4164_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4164_2), .COMP_OUT(1'b0) );
// C_////Bridge      x86y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4165_5 ( .OUT(na4165_2), .IN1(na3_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y63     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4166_5 ( .OUT(na4166_2), .IN1(na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x156y86     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4167_5 ( .OUT(na4167_2), .IN1(1'b0), .IN2(na12_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x158y80     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4168_5 ( .OUT(na4168_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na12_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4169_5 ( .OUT(na4169_2), .IN1(1'b0), .IN2(1'b0), .IN3(na15_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4170_5 ( .OUT(na4170_2), .IN1(na16_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4171_5 ( .OUT(na4171_2), .IN1(na21_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4172_5 ( .OUT(na4172_2), .IN1(na21_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y79     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4173_5 ( .OUT(na4173_2), .IN1(na21_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4174_5 ( .OUT(na4174_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na25_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4175_5 ( .OUT(na4175_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na25_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x130y79     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4176_5 ( .OUT(na4176_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na25_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y82     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4177_5 ( .OUT(na4177_2), .IN1(na26_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y90     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4178_5 ( .OUT(na4178_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na26_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y80     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4179_5 ( .OUT(na4179_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na218_1) );
// C_////Bridge      x84y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4180_5 ( .OUT(na4180_2), .IN1(1'b0), .IN2(na223_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4181_5 ( .OUT(na4181_2), .IN1(1'b0), .IN2(1'b0), .IN3(na225_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4182_5 ( .OUT(na4182_2), .IN1(na234_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y81     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4183_5 ( .OUT(na4183_2), .IN1(na234_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4184_5 ( .OUT(na4184_2), .IN1(na234_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y80     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4185_5 ( .OUT(na4185_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na239_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4186_5 ( .OUT(na4186_2), .IN1(1'b0), .IN2(na241_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y83     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4187_5 ( .OUT(na4187_2), .IN1(1'b0), .IN2(1'b0), .IN3(na242_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y82     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4188_5 ( .OUT(na4188_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na245_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y84     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4189_5 ( .OUT(na4189_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na248_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y88     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4190_5 ( .OUT(na4190_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na253_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x132y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4191_5 ( .OUT(na4191_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na264_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x129y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4192_5 ( .OUT(na4192_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na277_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4193_5 ( .OUT(na4193_2), .IN1(1'b0), .IN2(1'b0), .IN3(na295_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4194_5 ( .OUT(na4194_2), .IN1(1'b0), .IN2(1'b0), .IN3(na316_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4195_5 ( .OUT(na4195_2), .IN1(1'b0), .IN2(1'b0), .IN3(na316_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x141y81     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4196_5 ( .OUT(na4196_2), .IN1(1'b0), .IN2(1'b0), .IN3(na349_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4197_5 ( .OUT(na4197_2), .IN1(1'b0), .IN2(1'b0), .IN3(na353_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y59     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4198_5 ( .OUT(na4198_2), .IN1(1'b0), .IN2(na389_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x146y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4199_5 ( .OUT(na4199_2), .IN1(1'b0), .IN2(1'b0), .IN3(na458_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y61     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4200_5 ( .OUT(na4200_2), .IN1(na530_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y59     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4201_5 ( .OUT(na4201_2), .IN1(na530_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x142y63     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4202_5 ( .OUT(na4202_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na539_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y85     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4203_5 ( .OUT(na4203_2), .IN1(na556_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y84     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4204_5 ( .OUT(na4204_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na565_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4205_5 ( .OUT(na4205_2), .IN1(1'b0), .IN2(1'b0), .IN3(na566_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4206_5 ( .OUT(na4206_2), .IN1(1'b0), .IN2(1'b0), .IN3(na566_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4207_5 ( .OUT(na4207_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na567_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x129y96     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4208_5 ( .OUT(na4208_2), .IN1(na570_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y91     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4209_5 ( .OUT(na4209_2), .IN1(na570_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4210_5 ( .OUT(na4210_2), .IN1(na571_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y72     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4211_5 ( .OUT(na4211_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na574_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4212_5 ( .OUT(na4212_2), .IN1(na575_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4213_5 ( .OUT(na4213_2), .IN1(na576_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y85     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4214_5 ( .OUT(na4214_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na577_1), .IN8(1'b0) );
// C_////Bridge      x117y90     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4215_5 ( .OUT(na4215_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na578_1), .IN8(1'b0) );
// C_////Bridge      x106y83     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4216_5 ( .OUT(na4216_2), .IN1(na580_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y86     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4217_5 ( .OUT(na4217_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na581_1), .IN8(1'b0) );
// C_////Bridge      x101y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4218_5 ( .OUT(na4218_2), .IN1(1'b0), .IN2(1'b0), .IN3(na582_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4219_5 ( .OUT(na4219_2), .IN1(1'b0), .IN2(1'b0), .IN3(na582_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4220_5 ( .OUT(na4220_2), .IN1(1'b0), .IN2(na585_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4221_5 ( .OUT(na4221_2), .IN1(na592_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4222_5 ( .OUT(na4222_2), .IN1(1'b0), .IN2(1'b0), .IN3(na598_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4223_5 ( .OUT(na4223_2), .IN1(na599_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4224_5 ( .OUT(na4224_2), .IN1(na599_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y74     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4225_5 ( .OUT(na4225_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na603_1), .IN8(1'b0) );
// C_////Bridge      x121y91     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4226_5 ( .OUT(na4226_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na612_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y68     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4227_5 ( .OUT(na4227_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na615_1) );
// C_////Bridge      x108y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4228_5 ( .OUT(na4228_2), .IN1(na658_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y96     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4229_5 ( .OUT(na4229_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na674_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y90     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4230_5 ( .OUT(na4230_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na677_1) );
// C_////Bridge      x122y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4231_5 ( .OUT(na4231_2), .IN1(na746_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4232_5 ( .OUT(na4232_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na747_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y72     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4233_5 ( .OUT(na4233_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na749_1) );
// C_////Bridge      x100y63     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4234_5 ( .OUT(na4234_2), .IN1(na750_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x131y96     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4235_5 ( .OUT(na4235_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na761_1) );
// C_////Bridge      x132y95     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4236_5 ( .OUT(na4236_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na762_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4237_5 ( .OUT(na4237_2), .IN1(1'b0), .IN2(1'b0), .IN3(na769_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4238_5 ( .OUT(na4238_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na771_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y94     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4239_5 ( .OUT(na4239_2), .IN1(na773_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y98     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4240_5 ( .OUT(na4240_2), .IN1(1'b0), .IN2(1'b0), .IN3(na809_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y87     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4241_5 ( .OUT(na4241_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na818_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4242_5 ( .OUT(na4242_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na821_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4243_5 ( .OUT(na4243_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na821_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4244_5 ( .OUT(na4244_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na821_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4245_5 ( .OUT(na4245_2), .IN1(1'b0), .IN2(na822_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y101     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4246_5 ( .OUT(na4246_2), .IN1(1'b0), .IN2(1'b0), .IN3(na824_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4247_5 ( .OUT(na4247_2), .IN1(1'b0), .IN2(1'b0), .IN3(na824_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4248_5 ( .OUT(na4248_2), .IN1(1'b0), .IN2(na827_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4249_5 ( .OUT(na4249_2), .IN1(1'b0), .IN2(na827_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y104     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4250_5 ( .OUT(na4250_2), .IN1(1'b0), .IN2(na827_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4251_5 ( .OUT(na4251_2), .IN1(1'b0), .IN2(na827_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y92     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4252_5 ( .OUT(na4252_2), .IN1(1'b0), .IN2(na829_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y95     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4253_5 ( .OUT(na4253_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na836_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y93     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4254_5 ( .OUT(na4254_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na836_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y98     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4255_5 ( .OUT(na4255_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na842_2), .IN8(1'b0) );
// C_////Bridge      x91y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4256_5 ( .OUT(na4256_2), .IN1(1'b0), .IN2(na844_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4257_5 ( .OUT(na4257_2), .IN1(1'b0), .IN2(na844_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y95     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4258_5 ( .OUT(na4258_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na845_1) );
// C_////Bridge      x89y86     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4259_5 ( .OUT(na4259_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na849_1) );
// C_////Bridge      x86y99     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4260_5 ( .OUT(na4260_2), .IN1(na854_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4261_5 ( .OUT(na4261_2), .IN1(1'b0), .IN2(na865_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y90     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4262_5 ( .OUT(na4262_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na869_1) );
// C_////Bridge      x88y71     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4263_5 ( .OUT(na4263_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na875_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x152y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4264_5 ( .OUT(na4264_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na882_1) );
// C_////Bridge      x150y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4265_5 ( .OUT(na4265_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na889_1) );
// C_////Bridge      x148y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4266_5 ( .OUT(na4266_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na891_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4267_5 ( .OUT(na4267_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na894_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y95     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4268_5 ( .OUT(na4268_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na898_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y102     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4269_5 ( .OUT(na4269_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na899_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4270_5 ( .OUT(na4270_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na899_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x141y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4271_5 ( .OUT(na4271_2), .IN1(1'b0), .IN2(na900_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y98     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4272_5 ( .OUT(na4272_2), .IN1(1'b0), .IN2(na900_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y97     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4273_5 ( .OUT(na4273_2), .IN1(1'b0), .IN2(1'b0), .IN3(na901_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x143y96     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4274_5 ( .OUT(na4274_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na901_2), .IN8(1'b0) );
// C_////Bridge      x145y98     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4275_5 ( .OUT(na4275_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na903_2) );
// C_////Bridge      x158y101     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4276_5 ( .OUT(na4276_2), .IN1(na906_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y96     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4277_5 ( .OUT(na4277_2), .IN1(1'b0), .IN2(1'b0), .IN3(na921_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y96     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4278_5 ( .OUT(na4278_2), .IN1(1'b0), .IN2(1'b0), .IN3(na921_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y99     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4279_5 ( .OUT(na4279_2), .IN1(na927_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x152y95     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4280_5 ( .OUT(na4280_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na929_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y96     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4281_5 ( .OUT(na4281_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na932_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y100     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4282_5 ( .OUT(na4282_2), .IN1(1'b0), .IN2(na933_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x146y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4283_5 ( .OUT(na4283_2), .IN1(na934_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y100     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4284_5 ( .OUT(na4284_2), .IN1(1'b0), .IN2(na938_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y99     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4285_5 ( .OUT(na4285_2), .IN1(na940_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x152y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4286_5 ( .OUT(na4286_2), .IN1(1'b0), .IN2(na946_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y88     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4287_5 ( .OUT(na4287_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na965_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y98     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4288_5 ( .OUT(na4288_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na977_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4289_5 ( .OUT(na4289_2), .IN1(na977_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y100     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4290_5 ( .OUT(na4290_2), .IN1(na977_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y95     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4291_5 ( .OUT(na4291_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na978_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4292_5 ( .OUT(na4292_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na978_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4293_5 ( .OUT(na4293_2), .IN1(1'b0), .IN2(na979_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4294_5 ( .OUT(na4294_2), .IN1(1'b0), .IN2(na979_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y98     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4295_5 ( .OUT(na4295_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na981_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y98     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4296_5 ( .OUT(na4296_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na981_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4297_5 ( .OUT(na4297_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na981_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y102     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4298_5 ( .OUT(na4298_2), .IN1(1'b0), .IN2(na984_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4299_5 ( .OUT(na4299_2), .IN1(1'b0), .IN2(1'b0), .IN3(na996_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y99     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4300_5 ( .OUT(na4300_2), .IN1(na1002_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4301_5 ( .OUT(na4301_2), .IN1(na1003_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y100     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4302_5 ( .OUT(na4302_2), .IN1(na1003_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y104     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4303_5 ( .OUT(na4303_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1006_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y101     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4304_5 ( .OUT(na4304_2), .IN1(na1007_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y100     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4305_5 ( .OUT(na4305_2), .IN1(na1008_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4306_5 ( .OUT(na4306_2), .IN1(na1008_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4307_5 ( .OUT(na4307_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1013_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y103     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4308_5 ( .OUT(na4308_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1023_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4309_5 ( .OUT(na4309_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1030_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x154y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4310_5 ( .OUT(na4310_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1034_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4311_5 ( .OUT(na4311_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1035_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x154y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4312_5 ( .OUT(na4312_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1048_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x154y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4313_5 ( .OUT(na4313_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1050_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4314_5 ( .OUT(na4314_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1142_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x129y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4315_5 ( .OUT(na4315_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1142_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4316_5 ( .OUT(na4316_2), .IN1(1'b0), .IN2(na1151_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y88     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4317_5 ( .OUT(na4317_2), .IN1(1'b0), .IN2(na1151_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y93     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4318_5 ( .OUT(na4318_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1154_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y94     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4319_5 ( .OUT(na4319_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1156_1) );
// C_////Bridge      x90y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4320_5 ( .OUT(na4320_2), .IN1(1'b0), .IN2(na1166_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y97     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4321_5 ( .OUT(na4321_2), .IN1(na1168_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y99     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4322_5 ( .OUT(na4322_2), .IN1(na1170_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4323_5 ( .OUT(na4323_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1182_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y98     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4324_5 ( .OUT(na4324_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1182_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x155y101     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4325_5 ( .OUT(na4325_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1184_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4326_5 ( .OUT(na4326_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1198_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y95     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4327_5 ( .OUT(na4327_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1200_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4328_5 ( .OUT(na4328_2), .IN1(1'b0), .IN2(na1214_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x153y63     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4329_5 ( .OUT(na4329_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1217_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4330_5 ( .OUT(na4330_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1224_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y80     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4331_5 ( .OUT(na4331_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1235_1) );
// C_////Bridge      x153y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4332_5 ( .OUT(na4332_2), .IN1(na1236_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x155y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4333_5 ( .OUT(na4333_2), .IN1(na1236_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y69     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4334_5 ( .OUT(na4334_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1238_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x152y70     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4335_5 ( .OUT(na4335_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1243_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4336_5 ( .OUT(na4336_2), .IN1(na1245_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4337_5 ( .OUT(na4337_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1246_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x154y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4338_5 ( .OUT(na4338_2), .IN1(1'b0), .IN2(na1251_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x152y72     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4339_5 ( .OUT(na4339_2), .IN1(1'b0), .IN2(na1251_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x156y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4340_5 ( .OUT(na4340_2), .IN1(1'b0), .IN2(na1251_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4341_5 ( .OUT(na4341_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1335_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4342_5 ( .OUT(na4342_2), .IN1(na1335_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y68     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4343_5 ( .OUT(na4343_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1343_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y78     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4344_5 ( .OUT(na4344_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1343_2), .IN8(1'b0) );
// C_////Bridge      x149y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4345_5 ( .OUT(na4345_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1386_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y77     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4346_5 ( .OUT(na4346_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1389_1) );
// C_////Bridge      x116y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4347_5 ( .OUT(na4347_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1400_1) );
// C_////Bridge      x92y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4348_5 ( .OUT(na4348_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1419_1) );
// C_////Bridge      x137y78     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4349_5 ( .OUT(na4349_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1451_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x135y82     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4350_5 ( .OUT(na4350_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1451_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4351_5 ( .OUT(na4351_2), .IN1(1'b0), .IN2(na1464_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x130y74     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4352_5 ( .OUT(na4352_2), .IN1(1'b0), .IN2(na1464_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4353_5 ( .OUT(na4353_2), .IN1(1'b0), .IN2(na1482_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y59     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4354_5 ( .OUT(na4354_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1500_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x140y94     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4355_5 ( .OUT(na4355_2), .IN1(1'b0), .IN2(na1513_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y63     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4356_5 ( .OUT(na4356_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1516_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y62     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4357_5 ( .OUT(na4357_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1620_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y96     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4358_5 ( .OUT(na4358_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1624_2) );
// C_////Bridge      x109y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4359_5 ( .OUT(na4359_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1638_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y81     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4360_5 ( .OUT(na4360_2), .IN1(na1811_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4361_5 ( .OUT(na4361_2), .IN1(1'b0), .IN2(na1824_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y90     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4362_5 ( .OUT(na4362_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1842_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x157y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4363_5 ( .OUT(na4363_2), .IN1(1'b0), .IN2(na1847_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y102     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4364_5 ( .OUT(na4364_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1852_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y65     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4365_5 ( .OUT(na4365_2), .IN1(1'b0), .IN2(na1859_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4366_5 ( .OUT(na4366_2), .IN1(1'b0), .IN2(na1859_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y74     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4367_5 ( .OUT(na4367_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3196_2), .IN8(1'b0) );
// C_////Bridge      x86y58     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4368_5 ( .OUT(na4368_2), .IN1(na3223_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4369_5 ( .OUT(na4369_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3290_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4370_5 ( .OUT(na4370_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3298_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4371_5 ( .OUT(na4371_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3363_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4372_5 ( .OUT(na4372_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3368_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4373_5 ( .OUT(na4373_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3454_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y94     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4374_5 ( .OUT(na4374_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3456_2) );
// C_////Bridge      x87y96     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4375_5 ( .OUT(na4375_2), .IN1(na3457_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y95     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4376_5 ( .OUT(na4376_2), .IN1(na3457_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y98     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4377_5 ( .OUT(na4377_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3457_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y85     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4378_5 ( .OUT(na4378_2), .IN1(na3470_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4379_5 ( .OUT(na4379_2), .IN1(na3471_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y88     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4380_5 ( .OUT(na4380_2), .IN1(1'b0), .IN2(na3477_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y71     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4381_5 ( .OUT(na4381_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3555_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y81     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4382_5 ( .OUT(na4382_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3646_2) );
// C_////Bridge      x150y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4383_5 ( .OUT(na4383_2), .IN1(1'b0), .IN2(na3656_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4384_5 ( .OUT(na4384_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3662_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y92     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4385_5 ( .OUT(na4385_2), .IN1(na3706_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y100     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4386_5 ( .OUT(na4386_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3711_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y98     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4387_5 ( .OUT(na4387_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3723_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y97     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4388_5 ( .OUT(na4388_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3728_1) );
// C_////Bridge      x135y79     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4389_5 ( .OUT(na4389_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3730_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4390_5 ( .OUT(na4390_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3735_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y84     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4391_5 ( .OUT(na4391_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3736_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y74     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4392_5 ( .OUT(na4392_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3739_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4393_5 ( .OUT(na4393_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3740_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x132y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4394_5 ( .OUT(na4394_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3741_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4395_5 ( .OUT(na4395_2), .IN1(1'b0), .IN2(na3742_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x155y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4396_5 ( .OUT(na4396_2), .IN1(na3744_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x156y97     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4397_5 ( .OUT(na4397_2), .IN1(na3744_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x157y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4398_5 ( .OUT(na4398_2), .IN1(1'b0), .IN2(na3745_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y100     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4399_5 ( .OUT(na4399_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3753_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x151y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4400_5 ( .OUT(na4400_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3759_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x154y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4401_5 ( .OUT(na4401_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3759_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x147y99     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4402_5 ( .OUT(na4402_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3763_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x156y99     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4403_5 ( .OUT(na4403_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3765_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x141y100     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4404_5 ( .OUT(na4404_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3766_2), .IN8(1'b0) );
// C_////Bridge      x153y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4405_5 ( .OUT(na4405_2), .IN1(1'b0), .IN2(na3768_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x158y98     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4406_5 ( .OUT(na4406_2), .IN1(1'b0), .IN2(na3768_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x150y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4407_5 ( .OUT(na4407_2), .IN1(1'b0), .IN2(na3770_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y97     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4408_5 ( .OUT(na4408_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3775_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x152y91     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4409_5 ( .OUT(na4409_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3776_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y87     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4410_5 ( .OUT(na4410_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3779_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x148y88     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4411_5 ( .OUT(na4411_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3780_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x149y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4412_5 ( .OUT(na4412_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3781_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x145y79     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4413_5 ( .OUT(na4413_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3782_2) );
// C_////Bridge      x143y74     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4414_5 ( .OUT(na4414_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3783_1), .IN8(1'b0) );
// C_////Bridge      x98y95     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4415_5 ( .OUT(na4415_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3793_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4416_5 ( .OUT(na4416_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3793_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y100     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4417_5 ( .OUT(na4417_2), .IN1(na3798_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4418_5 ( .OUT(na4418_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3800_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4419_5 ( .OUT(na4419_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3800_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y103     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4420_5 ( .OUT(na4420_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3802_2) );
// C_////Bridge      x106y101     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4421_5 ( .OUT(na4421_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3804_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4422_5 ( .OUT(na4422_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3808_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y90     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4423_5 ( .OUT(na4423_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3809_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x142y90     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4424_5 ( .OUT(na4424_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3814_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x144y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4425_5 ( .OUT(na4425_2), .IN1(1'b0), .IN2(na3815_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x139y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4426_5 ( .OUT(na4426_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3818_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x138y87     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4427_5 ( .OUT(na4427_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3819_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x135y85     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4428_5 ( .OUT(na4428_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3820_1) );
// C_////Bridge      x142y77     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4429_5 ( .OUT(na4429_2), .IN1(1'b0), .IN2(na3821_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x137y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4430_5 ( .OUT(na4430_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3822_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y79     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4431_5 ( .OUT(na4431_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3871_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y92     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4432_5 ( .OUT(na4432_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na4106_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y68     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4433_5 ( .OUT(na4433_2), .IN1(1'b0), .IN2(1'b0), .IN3(na4155_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_CP_route////      x79y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4434_1 ( .OUT(na4434_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x80y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4435_1 ( .OUT(na4435_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x81y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4436_1 ( .OUT(na4436_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x82y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4437_1 ( .OUT(na4437_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x83y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4438_1 ( .OUT(na4438_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x84y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4439_1 ( .OUT(na4439_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x85y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4440_1 ( .OUT(na4440_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x86y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4441_1 ( .OUT(na4441_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x87y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4442_1 ( .OUT(na4442_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x88y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4443_1 ( .OUT(na4443_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x89y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4444_1 ( .OUT(na4444_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x90y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4445_1 ( .OUT(na4445_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x91y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4446_1 ( .OUT(na4446_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x92y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4447_1 ( .OUT(na4447_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x93y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4448_1 ( .OUT(na4448_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x94y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4449_1 ( .OUT(na4449_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x95y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4450_1 ( .OUT(na4450_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x96y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4451_1 ( .OUT(na4451_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x97y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4452_1 ( .OUT(na4452_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x98y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4453_1 ( .OUT(na4453_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x99y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4454_1 ( .OUT(na4454_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x100y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4455_1 ( .OUT(na4455_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x101y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4456_1 ( .OUT(na4456_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x102y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4457_1 ( .OUT(na4457_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x103y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4458_1 ( .OUT(na4458_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x104y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4459_1 ( .OUT(na4459_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x105y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4460_1 ( .OUT(na4460_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x106y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4461_1 ( .OUT(na4461_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x107y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4462_1 ( .OUT(na4462_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x108y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4463_1 ( .OUT(na4463_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x109y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4464_1 ( .OUT(na4464_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x110y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4465_1 ( .OUT(na4465_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x111y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4466_1 ( .OUT(na4466_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x112y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4467_1 ( .OUT(na4467_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x113y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4468_1 ( .OUT(na4468_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x114y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4469_1 ( .OUT(na4469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x115y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4470_1 ( .OUT(na4470_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x116y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4471_1 ( .OUT(na4471_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x117y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4472_1 ( .OUT(na4472_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x118y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4473_1 ( .OUT(na4473_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x119y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4474_1 ( .OUT(na4474_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x120y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4475_1 ( .OUT(na4475_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x121y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4476_1 ( .OUT(na4476_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x122y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4477_1 ( .OUT(na4477_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x123y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4478_1 ( .OUT(na4478_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x124y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4479_1 ( .OUT(na4479_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x125y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4480_1 ( .OUT(na4480_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x126y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4481_1 ( .OUT(na4481_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x127y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4482_1 ( .OUT(na4482_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x128y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4483_1 ( .OUT(na4483_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x129y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4484_1 ( .OUT(na4484_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x130y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4485_1 ( .OUT(na4485_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x131y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4486_1 ( .OUT(na4486_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x132y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4487_1 ( .OUT(na4487_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x133y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4488_1 ( .OUT(na4488_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x134y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4489_1 ( .OUT(na4489_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x135y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4490_1 ( .OUT(na4490_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x136y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4491_1 ( .OUT(na4491_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x137y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4492_1 ( .OUT(na4492_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x138y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4493_1 ( .OUT(na4493_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x139y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4494_1 ( .OUT(na4494_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x140y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4495_1 ( .OUT(na4495_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x141y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4496_1 ( .OUT(na4496_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x142y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4497_1 ( .OUT(na4497_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x143y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4498_1 ( .OUT(na4498_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x144y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4499_1 ( .OUT(na4499_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x145y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4500_1 ( .OUT(na4500_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x146y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4501_1 ( .OUT(na4501_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x147y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4502_1 ( .OUT(na4502_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x148y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4503_1 ( .OUT(na4503_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x149y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4504_1 ( .OUT(na4504_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x150y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4505_1 ( .OUT(na4505_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x151y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4506_1 ( .OUT(na4506_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x152y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4507_1 ( .OUT(na4507_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x153y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4508_1 ( .OUT(na4508_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x154y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4509_1 ( .OUT(na4509_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x155y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4510_1 ( .OUT(na4510_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x156y56     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a4511_1 ( .OUT(na4511_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x78y56     80'h00_0078_09_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4512_1 ( .OUT(na4512_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1923_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4512_4 ( .OUT(na4512_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na25_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9000)) 
           _a4512_6 ( .COUTX(na4512_3), .POUTX(na4512_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na4512_1), .OUT2(na4512_2), .COMP_OUT(1'b0) );
endmodule
