//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 Jul 2023)
//  Compile Time: 2023-07-20 13:23:25
//  Program Run:  2023-08-07 04:02:59
//  Program Call: ../../bin/p_r/p_r -i net/aes256_impl_synth.v -o aes256_impl -ccf src/aes256_impl.ccf 
//  File Type:    Verilog

// Gatecount:   1972
module aes256_impl (clk10 , reset_n ,
       led 
       ) ;

input  clk10;
input  reset_n;

output [7:0]led;



wire [7:0]led;
wire clk10;
wire na2_1;
wire na5_1;
wire na5_1_i;
wire na5_2;
wire na5_2_i;
wire na6_1;
wire na6_1_i;
wire na6_2;
wire na6_2_i;
wire na7_1;
wire na7_1_i;
wire na7_2;
wire na7_2_i;
wire na8_2;
wire na8_2_i;
wire na11_1;
wire na11_2;
wire na13_1;
wire na15_1;
wire na18_1;
wire na19_1;
wire na20_1;
wire na20_2;
wire na22_1;
wire na23_1;
wire na23_2;
wire na25_2;
wire na27_1;
wire na29_1;
wire na32_1;
wire na33_1;
wire na34_1;
wire na35_1;
wire na36_1;
wire na37_1;
wire na38_1;
wire na42_1;
wire na42_2;
wire na43_1;
wire na45_1;
wire na46_1;
wire na48_1;
wire na48_2;
wire na49_1;
wire na50_1;
wire na51_1;
wire na54_1;
wire na55_1;
wire na55_1_i;
wire na55_2;
wire na55_2_i;
wire na57_2;
wire na59_1;
wire na61_1;
wire na62_2;
wire na65_1;
wire na65_2;
wire na66_1;
wire na66_2;
wire na69_1;
wire na69_2;
wire na70_1;
wire na72_1;
wire na73_1;
wire na74_1;
wire na75_1;
wire na75_2;
wire na82_1;
wire na82_2;
wire na83_1;
wire na85_1;
wire na85_2;
wire na86_1;
wire na88_2;
wire na91_2;
wire na93_1;
wire na94_1;
wire na94_2;
wire na95_1;
wire na97_1;
wire na98_1;
wire na99_2;
wire na99_2_i;
wire na103_1;
wire na104_1;
wire na104_2;
wire na105_1;
wire na105_2;
wire na106_1;
wire na107_1;
wire na107_1_i;
wire na107_2;
wire na107_2_i;
wire na109_2;
wire na111_1;
wire na112_1;
wire na112_2;
wire na113_1;
wire na115_1;
wire na119_1;
wire na120_2;
wire na121_1;
wire na121_2;
wire na122_2;
wire na123_1;
wire na123_1_i;
wire na127_1;
wire na128_1;
wire na128_2;
wire na129_1;
wire na129_1_i;
wire na129_2;
wire na129_2_i;
wire na133_1;
wire na137_1;
wire na138_1;
wire na139_1;
wire na140_1;
wire na140_1_i;
wire na141_1;
wire na143_1;
wire na144_1;
wire na146_1;
wire na146_1_i;
wire na146_2;
wire na146_2_i;
wire na148_1;
wire na149_1;
wire na150_1;
wire na150_2;
wire na151_1;
wire na152_1;
wire na152_1_i;
wire na152_2;
wire na152_2_i;
wire na153_2;
wire na155_1;
wire na156_1;
wire na157_1;
wire na162_1;
wire na163_1;
wire na164_1;
wire na164_1_i;
wire na164_2;
wire na164_2_i;
wire na168_1;
wire na169_1;
wire na173_1;
wire na175_1;
wire na176_1;
wire na176_1_i;
wire na176_2;
wire na176_2_i;
wire na178_1;
wire na178_2;
wire na180_1;
wire na181_1;
wire na182_1;
wire na183_1;
wire na184_2;
wire na184_2_i;
wire na188_1;
wire na189_1;
wire na190_1;
wire na190_1_i;
wire na190_2;
wire na190_2_i;
wire na193_1;
wire na194_1;
wire na195_2;
wire na196_1;
wire na196_1_i;
wire na196_2;
wire na196_2_i;
wire na199_1;
wire na200_1;
wire na201_1;
wire na202_1;
wire na202_1_i;
wire na202_2;
wire na202_2_i;
wire na205_1;
wire na207_1;
wire na208_1;
wire na208_1_i;
wire na208_2;
wire na208_2_i;
wire na209_1;
wire na211_1;
wire na212_1;
wire na213_1;
wire na214_1;
wire na214_1_i;
wire na214_2;
wire na214_2_i;
wire na215_1;
wire na217_1;
wire na218_1;
wire na220_1;
wire na220_1_i;
wire na223_1;
wire na224_1;
wire na225_1;
wire na226_2;
wire na226_2_i;
wire na227_2;
wire na229_1;
wire na230_1;
wire na231_1;
wire na235_1;
wire na237_1;
wire na242_1;
wire na243_1;
wire na245_1;
wire na247_1;
wire na248_1;
wire na249_1;
wire na253_1;
wire na255_1;
wire na256_1;
wire na256_1_i;
wire na258_1;
wire na258_2;
wire na260_1;
wire na261_1;
wire na265_1;
wire na267_1;
wire na268_1;
wire na268_1_i;
wire na271_1;
wire na272_1;
wire na273_1;
wire na273_1_i;
wire na274_1;
wire na276_1;
wire na277_1;
wire na278_1;
wire na278_1_i;
wire na279_2;
wire na281_1;
wire na282_1;
wire na283_1;
wire na283_1_i;
wire na284_1;
wire na286_1;
wire na287_1;
wire na288_1;
wire na288_1_i;
wire na289_2;
wire na291_1;
wire na292_1;
wire na293_1;
wire na293_1_i;
wire na294_2;
wire na296_1;
wire na297_1;
wire na298_1;
wire na298_1_i;
wire na299_2;
wire na301_1;
wire na302_1;
wire na303_1;
wire na303_1_i;
wire na304_2;
wire na306_1;
wire na307_1;
wire na308_1;
wire na308_1_i;
wire na309_1;
wire na311_1;
wire na312_1;
wire na313_1;
wire na313_1_i;
wire na314_2;
wire na316_1;
wire na317_1;
wire na318_1;
wire na318_1_i;
wire na319_1;
wire na321_1;
wire na322_1;
wire na323_1;
wire na323_1_i;
wire na324_1;
wire na326_1;
wire na327_1;
wire na328_1;
wire na328_1_i;
wire na329_1;
wire na331_1;
wire na332_1;
wire na333_1;
wire na333_1_i;
wire na334_2;
wire na336_1;
wire na337_1;
wire na338_1;
wire na338_1_i;
wire na339_2;
wire na341_1;
wire na342_1;
wire na343_1;
wire na343_1_i;
wire na344_2;
wire na346_1;
wire na347_1;
wire na348_1;
wire na348_1_i;
wire na349_1;
wire na351_1;
wire na352_1;
wire na353_1;
wire na353_1_i;
wire na354_1;
wire na356_1;
wire na357_1;
wire na358_1;
wire na358_1_i;
wire na359_1;
wire na361_1;
wire na362_1;
wire na363_1;
wire na363_1_i;
wire na364_2;
wire na366_1;
wire na367_1;
wire na368_1;
wire na368_1_i;
wire na369_2;
wire na371_1;
wire na372_1;
wire na373_1;
wire na373_1_i;
wire na374_2;
wire na376_1;
wire na377_1;
wire na378_1;
wire na378_1_i;
wire na379_1;
wire na381_1;
wire na382_1;
wire na383_1;
wire na383_1_i;
wire na384_2;
wire na386_1;
wire na387_1;
wire na388_1;
wire na388_1_i;
wire na389_1;
wire na391_1;
wire na392_1;
wire na393_1;
wire na393_1_i;
wire na394_1;
wire na396_1;
wire na397_1;
wire na398_1;
wire na398_1_i;
wire na399_1;
wire na401_1;
wire na402_1;
wire na403_1;
wire na403_1_i;
wire na404_2;
wire na406_1;
wire na407_1;
wire na408_1;
wire na408_1_i;
wire na409_2;
wire na411_1;
wire na412_1;
wire na413_1;
wire na413_1_i;
wire na414_2;
wire na416_1;
wire na417_1;
wire na418_1;
wire na418_1_i;
wire na419_1;
wire na421_1;
wire na422_1;
wire na423_1;
wire na423_1_i;
wire na424_1;
wire na426_1;
wire na427_1;
wire na428_1;
wire na428_1_i;
wire na429_1;
wire na430_1;
wire na430_1_i;
wire na430_2;
wire na430_2_i;
wire na431_1;
wire na431_1_i;
wire na432_2;
wire na432_2_i;
wire na433_1;
wire na433_1_i;
wire na434_2;
wire na434_2_i;
wire na435_1;
wire na435_1_i;
wire na436_2;
wire na436_2_i;
wire na437_2;
wire na437_2_i;
wire na438_1;
wire na438_1_i;
wire na438_2;
wire na438_2_i;
wire na439_2;
wire na439_2_i;
wire na440_1;
wire na440_1_i;
wire na441_2;
wire na441_2_i;
wire na442_1;
wire na442_1_i;
wire na443_2;
wire na443_2_i;
wire na444_2;
wire na444_2_i;
wire na445_1;
wire na445_1_i;
wire na446_2;
wire na446_2_i;
wire na447_1;
wire na447_1_i;
wire na448_2;
wire na448_2_i;
wire na449_1;
wire na449_1_i;
wire na450_1;
wire na450_1_i;
wire na450_2;
wire na450_2_i;
wire na451_1;
wire na451_1_i;
wire na452_1;
wire na452_1_i;
wire na452_2;
wire na452_2_i;
wire na453_1;
wire na453_1_i;
wire na454_2;
wire na454_2_i;
wire na455_1;
wire na455_1_i;
wire na456_2;
wire na456_2_i;
wire na457_1;
wire na457_1_i;
wire na458_2;
wire na458_2_i;
wire na459_2;
wire na459_2_i;
wire na460_2;
wire na460_2_i;
wire na461_1;
wire na461_1_i;
wire na461_2;
wire na461_2_i;
wire na462_1;
wire na462_1_i;
wire na462_2;
wire na462_2_i;
wire na463_2;
wire na463_2_i;
wire na464_2;
wire na464_2_i;
wire na465_1;
wire na465_1_i;
wire na466_1;
wire na466_1_i;
wire na467_1;
wire na467_1_i;
wire na467_2;
wire na467_2_i;
wire na468_1;
wire na468_1_i;
wire na468_2;
wire na468_2_i;
wire na469_2;
wire na469_2_i;
wire na470_1;
wire na470_1_i;
wire na470_2;
wire na470_2_i;
wire na471_1;
wire na471_1_i;
wire na472_2;
wire na472_2_i;
wire na473_2;
wire na473_2_i;
wire na474_2;
wire na474_2_i;
wire na475_1;
wire na475_1_i;
wire na476_1;
wire na476_1_i;
wire na477_1;
wire na477_1_i;
wire na478_1;
wire na478_1_i;
wire na478_2;
wire na478_2_i;
wire na479_2;
wire na479_2_i;
wire na480_2;
wire na480_2_i;
wire na481_2;
wire na481_2_i;
wire na482_1;
wire na482_1_i;
wire na483_2;
wire na483_2_i;
wire na484_2;
wire na484_2_i;
wire na485_1;
wire na485_1_i;
wire na486_1;
wire na486_1_i;
wire na487_1;
wire na487_1_i;
wire na488_2;
wire na488_2_i;
wire na489_2;
wire na489_2_i;
wire na490_1;
wire na490_1_i;
wire na490_2;
wire na490_2_i;
wire na491_2;
wire na491_2_i;
wire na492_1;
wire na492_1_i;
wire na492_2;
wire na492_2_i;
wire na493_1;
wire na493_1_i;
wire na495_1;
wire na495_1_i;
wire na496_1;
wire na496_1_i;
wire na497_2;
wire na497_2_i;
wire na498_2;
wire na498_2_i;
wire na499_2;
wire na499_2_i;
wire na500_1;
wire na500_1_i;
wire na501_1;
wire na501_1_i;
wire na503_1;
wire na503_1_i;
wire na504_2;
wire na504_2_i;
wire na505_2;
wire na505_2_i;
wire na506_2;
wire na506_2_i;
wire na507_1;
wire na507_1_i;
wire na508_1;
wire na508_1_i;
wire na509_1;
wire na509_1_i;
wire na510_2;
wire na510_2_i;
wire na511_1;
wire na511_1_i;
wire na512_2;
wire na512_2_i;
wire na513_2;
wire na513_2_i;
wire na515_2;
wire na515_2_i;
wire na517_1;
wire na517_1_i;
wire na518_1;
wire na518_1_i;
wire na519_1;
wire na519_1_i;
wire na520_2;
wire na520_2_i;
wire na521_2;
wire na521_2_i;
wire na522_2;
wire na522_2_i;
wire na523_1;
wire na523_1_i;
wire na524_1;
wire na524_1_i;
wire na525_1;
wire na525_1_i;
wire na526_2;
wire na526_2_i;
wire na527_2;
wire na527_2_i;
wire na528_2;
wire na528_2_i;
wire na529_1;
wire na529_1_i;
wire na530_1;
wire na530_1_i;
wire na531_1;
wire na531_1_i;
wire na532_2;
wire na532_2_i;
wire na533_2;
wire na533_2_i;
wire na534_2;
wire na534_2_i;
wire na535_1;
wire na535_1_i;
wire na536_2;
wire na536_2_i;
wire na537_1;
wire na537_1_i;
wire na538_2;
wire na538_2_i;
wire na539_2;
wire na539_2_i;
wire na540_1;
wire na540_1_i;
wire na541_1;
wire na541_1_i;
wire na542_2;
wire na542_2_i;
wire na543_2;
wire na543_2_i;
wire na544_2;
wire na544_2_i;
wire na545_1;
wire na545_1_i;
wire na546_1;
wire na546_1_i;
wire na547_1;
wire na547_1_i;
wire na548_2;
wire na548_2_i;
wire na549_2;
wire na549_2_i;
wire na550_2;
wire na550_2_i;
wire na551_1;
wire na551_1_i;
wire na552_1;
wire na552_1_i;
wire na553_1;
wire na553_1_i;
wire na554_2;
wire na554_2_i;
wire na555_2;
wire na555_2_i;
wire na556_2;
wire na556_2_i;
wire na557_1;
wire na557_1_i;
wire na558_2;
wire na558_2_i;
wire na559_1;
wire na559_1_i;
wire na560_1;
wire na560_1_i;
wire na561_1;
wire na561_1_i;
wire na562_2;
wire na562_2_i;
wire na563_2;
wire na563_2_i;
wire na564_2;
wire na564_2_i;
wire na565_1;
wire na565_1_i;
wire na566_1;
wire na566_1_i;
wire na567_1;
wire na567_1_i;
wire na568_1;
wire na568_1_i;
wire na569_1;
wire na569_1_i;
wire na570_1;
wire na570_1_i;
wire na571_1;
wire na571_1_i;
wire na572_2;
wire na572_2_i;
wire na573_1;
wire na573_1_i;
wire na574_2;
wire na574_2_i;
wire na575_1;
wire na575_1_i;
wire na576_2;
wire na576_2_i;
wire na577_1;
wire na577_1_i;
wire na578_2;
wire na578_2_i;
wire na579_1;
wire na579_1_i;
wire na580_2;
wire na580_2_i;
wire na581_1;
wire na581_1_i;
wire na582_2;
wire na582_2_i;
wire na583_1;
wire na583_1_i;
wire na584_2;
wire na584_2_i;
wire na585_1;
wire na585_1_i;
wire na586_2;
wire na586_2_i;
wire na587_1;
wire na587_1_i;
wire na588_2;
wire na588_2_i;
wire na589_1;
wire na589_1_i;
wire na591_2;
wire na591_2_i;
wire na592_1;
wire na592_1_i;
wire na593_2;
wire na593_2_i;
wire na594_1;
wire na594_1_i;
wire na595_2;
wire na595_2_i;
wire na596_1;
wire na596_1_i;
wire na597_2;
wire na597_2_i;
wire na599_1;
wire na599_1_i;
wire na600_2;
wire na600_2_i;
wire na601_1;
wire na601_1_i;
wire na602_2;
wire na602_2_i;
wire na603_1;
wire na603_1_i;
wire na604_2;
wire na604_2_i;
wire na605_1;
wire na605_1_i;
wire na606_2;
wire na606_2_i;
wire na607_1;
wire na607_1_i;
wire na608_2;
wire na608_2_i;
wire na609_1;
wire na609_1_i;
wire na611_2;
wire na611_2_i;
wire na615_1;
wire na615_1_i;
wire na616_2;
wire na616_2_i;
wire na617_1;
wire na617_1_i;
wire na618_2;
wire na618_2_i;
wire na621_1;
wire na621_1_i;
wire na622_2;
wire na622_2_i;
wire na623_1;
wire na623_1_i;
wire na624_2;
wire na624_2_i;
wire na625_2;
wire na625_2_i;
wire na626_2;
wire na626_2_i;
wire na627_1;
wire na627_1_i;
wire na628_1;
wire na628_1_i;
wire na629_2;
wire na629_2_i;
wire na630_1;
wire na630_1_i;
wire na631_1;
wire na631_1_i;
wire na632_1;
wire na632_1_i;
wire na633_2;
wire na633_2_i;
wire na634_1;
wire na634_1_i;
wire na635_2;
wire na635_2_i;
wire na636_1;
wire na636_1_i;
wire na637_2;
wire na637_2_i;
wire na638_1;
wire na638_1_i;
wire na639_2;
wire na639_2_i;
wire na640_1;
wire na640_1_i;
wire na641_2;
wire na641_2_i;
wire na642_1;
wire na642_1_i;
wire na643_2;
wire na643_2_i;
wire na644_1;
wire na644_1_i;
wire na645_2;
wire na645_2_i;
wire na646_1;
wire na646_1_i;
wire na647_2;
wire na647_2_i;
wire na648_1;
wire na648_1_i;
wire na649_2;
wire na649_2_i;
wire na650_1;
wire na650_1_i;
wire na651_2;
wire na651_2_i;
wire na652_1;
wire na652_1_i;
wire na653_2;
wire na653_2_i;
wire na654_1;
wire na654_1_i;
wire na655_2;
wire na655_2_i;
wire na656_1;
wire na656_1_i;
wire na657_2;
wire na657_2_i;
wire na658_1;
wire na658_1_i;
wire na659_2;
wire na659_2_i;
wire na660_1;
wire na660_1_i;
wire na661_2;
wire na661_2_i;
wire na662_1;
wire na662_1_i;
wire na663_2;
wire na663_2_i;
wire na664_1;
wire na664_1_i;
wire na665_2;
wire na665_2_i;
wire na666_1;
wire na666_1_i;
wire na667_2;
wire na667_2_i;
wire na668_1;
wire na668_1_i;
wire na669_2;
wire na669_2_i;
wire na670_1;
wire na670_1_i;
wire na671_2;
wire na671_2_i;
wire na672_1;
wire na672_1_i;
wire na673_2;
wire na673_2_i;
wire na674_1;
wire na674_1_i;
wire na675_2;
wire na675_2_i;
wire na676_1;
wire na676_1_i;
wire na677_2;
wire na677_2_i;
wire na678_1;
wire na678_1_i;
wire na679_2;
wire na679_2_i;
wire na680_1;
wire na680_1_i;
wire na681_2;
wire na681_2_i;
wire na682_1;
wire na682_1_i;
wire na683_2;
wire na683_2_i;
wire na684_1;
wire na684_1_i;
wire na685_1;
wire na685_1_i;
wire na685_2;
wire na685_2_i;
wire na686_1;
wire na686_2;
wire na688_1;
wire na688_1_i;
wire na688_2;
wire na688_2_i;
wire na690_1;
wire na690_1_i;
wire na690_2;
wire na690_2_i;
wire na692_2;
wire na692_2_i;
wire na693_1;
wire na693_2;
wire na695_2;
wire na696_1;
wire na697_1;
wire na699_1;
wire na700_1;
wire na700_2;
wire na702_1;
wire na702_2;
wire na703_1;
wire na703_2;
wire na704_1;
wire na704_2;
wire na706_1;
wire na706_2;
wire na707_1;
wire na709_1;
wire na711_1;
wire na713_1;
wire na716_1;
wire na717_1;
wire na718_1;
wire na719_1;
wire na720_1;
wire na721_1;
wire na722_1;
wire na723_1;
wire na724_1;
wire na725_2;
wire na726_1;
wire na727_1;
wire na729_1;
wire na729_2;
wire na730_1;
wire na732_1;
wire na733_1;
wire na734_1;
wire na735_1;
wire na736_1;
wire na737_1;
wire na738_1;
wire na738_1_i;
wire na739_1;
wire na739_2;
wire na741_2;
wire na742_1;
wire na743_1;
wire na744_1;
wire na746_1;
wire na747_1;
wire na747_1_i;
wire na748_1;
wire na748_2;
wire na749_1;
wire na750_1;
wire na752_2;
wire na753_1;
wire na753_1_i;
wire na754_1;
wire na754_2;
wire na755_1;
wire na757_1;
wire na758_1;
wire na759_1;
wire na759_1_i;
wire na760_1;
wire na760_2;
wire na761_1;
wire na763_1;
wire na763_1_i;
wire na764_1;
wire na764_2;
wire na765_1;
wire na766_1;
wire na768_1;
wire na768_1_i;
wire na769_1;
wire na769_2;
wire na770_1;
wire na770_1_i;
wire na771_1;
wire na771_2;
wire na772_2;
wire na773_1;
wire na773_1_i;
wire na774_1;
wire na774_2;
wire na775_1;
wire na776_2;
wire na777_1;
wire na778_1;
wire na779_1;
wire na780_2;
wire na781_1;
wire na781_2;
wire na783_1;
wire na783_2;
wire na784_1;
wire na786_1;
wire na789_1;
wire na791_1;
wire na794_1;
wire na795_2;
wire na796_1;
wire na797_1;
wire na800_1;
wire na801_1;
wire na802_1;
wire na803_1;
wire na804_1;
wire na806_1;
wire na807_2;
wire na808_1;
wire na809_1;
wire na810_1;
wire na811_1;
wire na812_1;
wire na814_1;
wire na815_1;
wire na816_2;
wire na817_1;
wire na818_1;
wire na819_1;
wire na819_1_i;
wire na820_1;
wire na820_2;
wire na821_1;
wire na822_1;
wire na823_1;
wire na824_1;
wire na825_1;
wire na826_1;
wire na827_1;
wire na828_1;
wire na828_1_i;
wire na829_1;
wire na829_2;
wire na830_2;
wire na831_1;
wire na832_1;
wire na832_1_i;
wire na833_1;
wire na833_2;
wire na834_2;
wire na836_1;
wire na837_1;
wire na838_1;
wire na838_1_i;
wire na839_1;
wire na839_2;
wire na840_1;
wire na841_1;
wire na841_1_i;
wire na842_1;
wire na842_2;
wire na844_1;
wire na844_1_i;
wire na845_1;
wire na845_2;
wire na846_1;
wire na846_1_i;
wire na847_1;
wire na847_2;
wire na848_1;
wire na848_1_i;
wire na849_1;
wire na849_2;
wire na850_1;
wire na851_1;
wire na851_2;
wire na852_1;
wire na853_1;
wire na856_1;
wire na858_1;
wire na858_2;
wire na860_1;
wire na860_2;
wire na862_1;
wire na863_1;
wire na865_1;
wire na868_1;
wire na869_1;
wire na870_2;
wire na874_1;
wire na875_1;
wire na876_1;
wire na877_1;
wire na878_1;
wire na878_2;
wire na879_2;
wire na880_1;
wire na881_1;
wire na882_1;
wire na883_1;
wire na884_1;
wire na888_1;
wire na889_1;
wire na890_1;
wire na891_1;
wire na892_1;
wire na894_1;
wire na895_2;
wire na896_1;
wire na897_1;
wire na898_1;
wire na898_1_i;
wire na899_1;
wire na899_2;
wire na900_1;
wire na900_2;
wire na901_1;
wire na904_1;
wire na905_1;
wire na906_1;
wire na907_1;
wire na907_1_i;
wire na908_1;
wire na908_2;
wire na911_1;
wire na911_1_i;
wire na912_1;
wire na912_2;
wire na913_1;
wire na915_1;
wire na916_1;
wire na917_1;
wire na917_1_i;
wire na918_1;
wire na918_2;
wire na919_2;
wire na920_1;
wire na920_1_i;
wire na921_1;
wire na921_2;
wire na923_1;
wire na924_1;
wire na924_1_i;
wire na925_1;
wire na925_2;
wire na926_1;
wire na926_1_i;
wire na927_1;
wire na927_2;
wire na928_1;
wire na928_1_i;
wire na929_1;
wire na929_1_i;
wire na930_1;
wire na930_1_i;
wire na931_1;
wire na931_1_i;
wire na932_1;
wire na932_1_i;
wire na933_1;
wire na933_1_i;
wire na934_1;
wire na934_1_i;
wire na935_1;
wire na935_1_i;
wire na936_1;
wire na936_1_i;
wire na937_1;
wire na937_1_i;
wire na938_1;
wire na938_1_i;
wire na939_1;
wire na939_1_i;
wire na940_1;
wire na940_1_i;
wire na941_1;
wire na941_1_i;
wire na942_1;
wire na942_1_i;
wire na943_1;
wire na943_1_i;
wire na944_1;
wire na944_1_i;
wire na945_1;
wire na945_1_i;
wire na946_1;
wire na946_1_i;
wire na947_1;
wire na947_1_i;
wire na948_1;
wire na948_1_i;
wire na949_1;
wire na949_1_i;
wire na950_1;
wire na950_1_i;
wire na951_1;
wire na951_1_i;
wire na952_1;
wire na952_1_i;
wire na953_1;
wire na953_1_i;
wire na954_1;
wire na954_1_i;
wire na955_1;
wire na955_1_i;
wire na956_1;
wire na956_1_i;
wire na957_1;
wire na957_1_i;
wire na958_1;
wire na958_1_i;
wire na959_1;
wire na959_1_i;
wire na960_1;
wire na960_1_i;
wire na961_1;
wire na961_1_i;
wire na962_1;
wire na962_1_i;
wire na963_1;
wire na963_1_i;
wire na964_1;
wire na964_1_i;
wire na965_1;
wire na965_1_i;
wire na966_1;
wire na966_1_i;
wire na967_1;
wire na967_1_i;
wire na968_1;
wire na968_1_i;
wire na969_1;
wire na969_1_i;
wire na970_1;
wire na970_1_i;
wire na971_1;
wire na971_1_i;
wire na972_1;
wire na972_1_i;
wire na973_1;
wire na973_1_i;
wire na974_1;
wire na974_1_i;
wire na975_1;
wire na975_1_i;
wire na976_1;
wire na976_1_i;
wire na977_1;
wire na977_1_i;
wire na978_1;
wire na978_1_i;
wire na979_1;
wire na979_1_i;
wire na980_1;
wire na980_1_i;
wire na981_1;
wire na981_1_i;
wire na982_1;
wire na982_1_i;
wire na983_1;
wire na983_1_i;
wire na984_1;
wire na984_1_i;
wire na985_1;
wire na985_1_i;
wire na986_1;
wire na986_1_i;
wire na987_1;
wire na987_1_i;
wire na988_1;
wire na988_1_i;
wire na989_1;
wire na989_1_i;
wire na990_1;
wire na990_1_i;
wire na991_1;
wire na991_1_i;
wire na992_1;
wire na992_1_i;
wire na993_1;
wire na993_1_i;
wire na994_1;
wire na994_1_i;
wire na995_1;
wire na995_1_i;
wire na996_1;
wire na996_1_i;
wire na997_1;
wire na997_1_i;
wire na998_1;
wire na998_1_i;
wire na999_1;
wire na999_1_i;
wire reset_n;
wire na1000_1;
wire na1000_1_i;
wire na1001_1;
wire na1001_1_i;
wire na1002_1;
wire na1002_1_i;
wire na1003_1;
wire na1003_1_i;
wire na1004_1;
wire na1004_1_i;
wire na1005_1;
wire na1005_1_i;
wire na1006_1;
wire na1006_1_i;
wire na1007_1;
wire na1007_1_i;
wire na1008_1;
wire na1008_1_i;
wire na1009_1;
wire na1009_2;
wire na1010_1;
wire na1010_2;
wire na1011_1;
wire na1011_2;
wire na1012_1;
wire na1012_2;
wire na1013_1;
wire na1013_2;
wire na1014_1;
wire na1014_2;
wire na1015_1;
wire na1015_2;
wire na1016_1;
wire na1016_2;
wire na1017_1;
wire na1017_2;
wire na1018_1;
wire na1018_1_i;
wire na1020_1;
wire na1021_1;
wire na1021_1_i;
wire na1022_1;
wire na1023_1;
wire na1023_1_i;
wire na1024_1;
wire na1025_1;
wire na1025_1_i;
wire na1026_1;
wire na1027_1;
wire na1027_1_i;
wire na1028_1;
wire na1029_1;
wire na1029_1_i;
wire na1030_1;
wire na1031_1;
wire na1031_1_i;
wire na1032_1;
wire na1033_1;
wire na1033_1_i;
wire na1034_1;
wire na1035_1;
wire na1035_1_i;
wire na1036_1;
wire na1037_1;
wire na1037_1_i;
wire na1038_1;
wire na1039_1;
wire na1039_1_i;
wire na1040_1;
wire na1041_1;
wire na1041_1_i;
wire na1042_1;
wire na1043_1;
wire na1043_1_i;
wire na1044_1;
wire na1045_1;
wire na1045_1_i;
wire na1046_1;
wire na1047_1;
wire na1047_1_i;
wire na1048_1;
wire na1049_1;
wire na1049_1_i;
wire na1050_1;
wire na1051_1;
wire na1051_1_i;
wire na1052_1;
wire na1053_1;
wire na1053_1_i;
wire na1054_1;
wire na1055_1;
wire na1055_1_i;
wire na1056_1;
wire na1057_1;
wire na1057_1_i;
wire na1058_1;
wire na1059_1;
wire na1059_1_i;
wire na1060_1;
wire na1061_1;
wire na1061_1_i;
wire na1062_1;
wire na1063_1;
wire na1063_1_i;
wire na1064_1;
wire na1065_1;
wire na1065_1_i;
wire na1066_1;
wire na1067_1;
wire na1067_1_i;
wire na1068_1;
wire na1069_1;
wire na1069_1_i;
wire na1070_1;
wire na1071_1;
wire na1071_1_i;
wire na1072_1;
wire na1073_1;
wire na1073_1_i;
wire na1074_1;
wire na1075_1;
wire na1075_1_i;
wire na1076_1;
wire na1077_1;
wire na1077_1_i;
wire na1078_1;
wire na1079_1;
wire na1079_1_i;
wire na1080_1;
wire na1081_1;
wire na1081_1_i;
wire na1082_1;
wire na1083_1;
wire na1083_1_i;
wire na1084_1;
wire na1084_1_i;
wire na1085_1;
wire na1085_1_i;
wire na1086_1;
wire na1087_1;
wire na1087_2;
wire na1089_1;
wire na1089_1_i;
wire na1089_2;
wire na1089_2_i;
wire na1090_2;
wire na1090_2_i;
wire na1091_1;
wire na1092_2;
wire na1094_1;
wire na1095_1;
wire na1096_1;
wire na1098_2;
wire na1099_2;
wire na1100_1;
wire na1101_1;
wire na1102_2;
wire na1103_1;
wire na1103_2;
wire na1104_1;
wire na1105_1;
wire na1106_1;
wire na1107_2;
wire na1108_1;
wire na1109_1;
wire na1110_1;
wire na1111_1;
wire na1112_1;
wire na1113_1;
wire na1114_1;
wire na1114_1_i;
wire na1115_1;
wire na1115_2;
wire na1116_1;
wire na1116_1_i;
wire na1117_2;
wire na1117_2_i;
wire na1118_2;
wire na1118_2_i;
wire na1120_1;
wire na1120_2;
wire na1121_1;
wire na1121_2;
wire na1122_2;
wire na1122_2_i;
wire na1123_1;
wire na1123_1_i;
wire na1124_1;
wire na1124_2;
wire na1125_2;
wire na1125_2_i;
wire na1126_1;
wire na1126_2;
wire na1127_1;
wire na1127_2;
wire na1128_1;
wire na1128_2;
wire na1129_1;
wire na1129_2;
wire na1130_1;
wire na1130_2;
wire na1131_1;
wire na1131_1_i;
wire na1132_1;
wire na1132_2;
wire na1133_2;
wire na1133_2_i;
wire na1134_1;
wire na1134_2;
wire na1135_1;
wire na1135_2;
wire na1136_1;
wire na1136_2;
wire na1137_1;
wire na1137_1_i;
wire na1138_2;
wire na1138_2_i;
wire na1139_1;
wire na1139_1_i;
wire na1140_1;
wire na1140_2;
wire na1141_1;
wire na1141_2;
wire na1142_2;
wire na1142_2_i;
wire na1143_1;
wire na1143_2;
wire na1144_1;
wire na1144_1_i;
wire na1145_2;
wire na1145_2_i;
wire na1146_1;
wire na1146_2;
wire na1147_1;
wire na1147_1_i;
wire na1148_2;
wire na1148_2_i;
wire na1149_1;
wire na1149_1_i;
wire na1150_1;
wire na1150_1_i;
wire na1151_2;
wire na1151_2_i;
wire na1152_1;
wire na1152_1_i;
wire na1153_2;
wire na1153_2_i;
wire na1154_1;
wire na1154_1_i;
wire na1155_1;
wire na1155_2;
wire na1156_2;
wire na1156_2_i;
wire na1157_2;
wire na1157_2_i;
wire na1158_1;
wire na1158_1_i;
wire na1159_2;
wire na1159_2_i;
wire na1160_1;
wire na1160_1_i;
wire na1161_1;
wire na1161_2;
wire na1162_1;
wire na1162_2;
wire na1163_1;
wire na1163_2;
wire na1164_2;
wire na1164_2_i;
wire na1165_1;
wire na1165_1_i;
wire na1166_1;
wire na1166_2;
wire na1167_2;
wire na1167_2_i;
wire na1168_1;
wire na1168_2;
wire na1169_2;
wire na1169_2_i;
wire na1170_1;
wire na1170_1_i;
wire na1171_1;
wire na1171_1_i;
wire na1172_2;
wire na1172_2_i;
wire na1173_1;
wire na1173_2;
wire na1174_1;
wire na1174_2;
wire na1175_1;
wire na1175_2;
wire na1176_1;
wire na1176_1_i;
wire na1177_2;
wire na1177_2_i;
wire na1178_1;
wire na1178_2;
wire na1179_1;
wire na1179_2;
wire na1180_1;
wire na1180_1_i;
wire na1181_2;
wire na1181_2_i;
wire na1182_1;
wire na1182_1_i;
wire na1183_1;
wire na1183_1_i;
wire na1184_1;
wire na1184_1_i;
wire na1185_1;
wire na1185_1_i;
wire na1186_2;
wire na1186_2_i;
wire na1187_1;
wire na1187_1_i;
wire na1188_2;
wire na1188_2_i;
wire na1189_1;
wire na1189_1_i;
wire na1190_2;
wire na1190_2_i;
wire na1191_1;
wire na1191_1_i;
wire na1192_1;
wire na1192_1_i;
wire na1193_2;
wire na1193_2_i;
wire na1194_1;
wire na1194_1_i;
wire na1195_2;
wire na1195_2_i;
wire na1196_2;
wire na1196_2_i;
wire na1197_2;
wire na1197_2_i;
wire na1198_1;
wire na1198_1_i;
wire na1199_1;
wire na1199_1_i;
wire na1200_2;
wire na1200_2_i;
wire na1201_2;
wire na1201_2_i;
wire na1202_1;
wire na1202_1_i;
wire na1203_1;
wire na1203_1_i;
wire na1204_2;
wire na1204_2_i;
wire na1205_1;
wire na1205_1_i;
wire na1206_2;
wire na1206_2_i;
wire na1207_1;
wire na1207_1_i;
wire na1208_2;
wire na1208_2_i;
wire na1209_2;
wire na1209_2_i;
wire na1210_2;
wire na1210_2_i;
wire na1211_1;
wire na1211_1_i;
wire na1212_2;
wire na1212_2_i;
wire na1213_1;
wire na1213_1_i;
wire na1214_1;
wire na1214_1_i;
wire na1215_1;
wire na1215_1_i;
wire na1216_1;
wire na1216_1_i;
wire na1217_2;
wire na1217_2_i;
wire na1218_1;
wire na1218_1_i;
wire na1219_1;
wire na1219_1_i;
wire na1220_2;
wire na1220_2_i;
wire na1221_1;
wire na1221_1_i;
wire na1222_1;
wire na1222_1_i;
wire na1223_2;
wire na1223_2_i;
wire na1224_2;
wire na1224_2_i;
wire na1225_2;
wire na1225_2_i;
wire na1226_1;
wire na1226_1_i;
wire na1227_1;
wire na1227_1_i;
wire na1228_2;
wire na1228_2_i;
wire na1229_1;
wire na1229_1_i;
wire na1230_1;
wire na1230_1_i;
wire na1231_2;
wire na1231_2_i;
wire na1232_2;
wire na1232_2_i;
wire na1233_1;
wire na1233_1_i;
wire na1234_1;
wire na1234_1_i;
wire na1235_1;
wire na1235_1_i;
wire na1236_2;
wire na1236_2_i;
wire na1237_1;
wire na1237_1_i;
wire na1238_1;
wire na1238_1_i;
wire na1239_1;
wire na1239_1_i;
wire na1240_1;
wire na1240_1_i;
wire na1241_1;
wire na1241_1_i;
wire na1242_2;
wire na1242_2_i;
wire na1243_1;
wire na1243_1_i;
wire na1244_1;
wire na1244_2;
wire na1245_2;
wire na1245_2_i;
wire na1246_1;
wire na1246_2;
wire na1247_1;
wire na1247_2;
wire na1248_1;
wire na1248_2;
wire na1249_1;
wire na1249_2;
wire na1250_1;
wire na1250_2;
wire na1251_1;
wire na1251_1_i;
wire na1252_1;
wire na1252_2;
wire na1253_2;
wire na1253_2_i;
wire na1254_1;
wire na1254_2;
wire na1255_1;
wire na1255_2;
wire na1256_1;
wire na1256_2;
wire na1257_1;
wire na1257_1_i;
wire na1258_2;
wire na1258_2_i;
wire na1259_1;
wire na1259_1_i;
wire na1260_1;
wire na1260_2;
wire na1261_1;
wire na1261_2;
wire na1262_2;
wire na1262_2_i;
wire na1263_1;
wire na1263_2;
wire na1264_1;
wire na1264_1_i;
wire na1265_2;
wire na1265_2_i;
wire na1266_1;
wire na1266_2;
wire na1267_1;
wire na1267_1_i;
wire na1268_2;
wire na1268_2_i;
wire na1269_1;
wire na1269_1_i;
wire na1270_1;
wire na1270_2;
wire na1271_1;
wire na1271_2;
wire na1272_2;
wire na1272_2_i;
wire na1273_1;
wire na1273_2;
wire na1274_1;
wire na1274_1_i;
wire na1275_2;
wire na1275_2_i;
wire na1276_1;
wire na1276_1_i;
wire na1277_2;
wire na1277_2_i;
wire na1278_2;
wire na1278_2_i;
wire na1279_1;
wire na1279_1_i;
wire na1280_2;
wire na1280_2_i;
wire na1281_1;
wire na1281_1_i;
wire na1282_2;
wire na1282_2_i;
wire na1283_1;
wire na1283_2;
wire na1284_1;
wire na1284_1_i;
wire na1285_2;
wire na1285_2_i;
wire na1286_2;
wire na1286_2_i;
wire na1287_1;
wire na1287_1_i;
wire na1288_2;
wire na1288_2_i;
wire na1289_1;
wire na1289_2;
wire na1290_1;
wire na1290_2;
wire na1291_1;
wire na1291_2;
wire na1292_1;
wire na1292_1_i;
wire na1293_2;
wire na1293_2_i;
wire na1294_1;
wire na1294_2;
wire na1295_1;
wire na1295_1_i;
wire na1296_1;
wire na1296_2;
wire na1297_1;
wire na1297_1_i;
wire na1298_2;
wire na1298_2_i;
wire na1299_2;
wire na1299_2_i;
wire na1300_1;
wire na1300_1_i;
wire na1301_2;
wire na1301_2_i;
wire na1302_1;
wire na1302_1_i;
wire na1303_2;
wire na1303_2_i;
wire na1304_1;
wire na1304_2;
wire na1305_1;
wire na1305_1_i;
wire na1306_1;
wire na1306_1_i;
wire na1307_2;
wire na1307_2_i;
wire na1308_1;
wire na1308_1_i;
wire na1309_1;
wire na1309_1_i;
wire na1310_1;
wire na1310_1_i;
wire na1311_2;
wire na1311_2_i;
wire na1312_2;
wire na1312_2_i;
wire na1313_1;
wire na1313_1_i;
wire na1314_1;
wire na1314_1_i;
wire na1315_2;
wire na1315_2_i;
wire na1316_1;
wire na1316_1_i;
wire na1317_2;
wire na1317_2_i;
wire na1318_1;
wire na1318_1_i;
wire na1319_2;
wire na1319_2_i;
wire na1320_2;
wire na1320_2_i;
wire na1321_1;
wire na1321_1_i;
wire na1322_2;
wire na1322_2_i;
wire na1323_1;
wire na1323_1_i;
wire na1324_2;
wire na1324_2_i;
wire na1325_2;
wire na1325_2_i;
wire na1326_2;
wire na1326_2_i;
wire na1327_2;
wire na1327_2_i;
wire na1328_1;
wire na1328_1_i;
wire na1329_1;
wire na1329_1_i;
wire na1330_1;
wire na1330_1_i;
wire na1331_2;
wire na1331_2_i;
wire na1332_2;
wire na1332_2_i;
wire na1333_1;
wire na1333_1_i;
wire na1334_1;
wire na1334_1_i;
wire na1335_1;
wire na1335_1_i;
wire na1336_2;
wire na1336_2_i;
wire na1337_2;
wire na1337_2_i;
wire na1338_2;
wire na1338_2_i;
wire na1339_2;
wire na1339_2_i;
wire na1340_1;
wire na1340_1_i;
wire na1341_1;
wire na1341_1_i;
wire na1342_2;
wire na1342_2_i;
wire na1343_1;
wire na1343_1_i;
wire na1344_2;
wire na1344_2_i;
wire na1345_1;
wire na1345_1_i;
wire na1346_2;
wire na1346_2_i;
wire na1347_2;
wire na1347_2_i;
wire na1348_1;
wire na1348_1_i;
wire na1349_1;
wire na1349_1_i;
wire na1350_2;
wire na1350_2_i;
wire na1351_1;
wire na1351_1_i;
wire na1352_2;
wire na1352_2_i;
wire na1353_1;
wire na1353_1_i;
wire na1354_2;
wire na1354_2_i;
wire na1355_2;
wire na1355_2_i;
wire na1356_1;
wire na1356_1_i;
wire na1357_2;
wire na1357_2_i;
wire na1358_2;
wire na1358_2_i;
wire na1359_1;
wire na1359_1_i;
wire na1360_2;
wire na1360_2_i;
wire na1361_1;
wire na1361_1_i;
wire na1362_2;
wire na1362_2_i;
wire na1363_1;
wire na1363_1_i;
wire na1364_1;
wire na1364_1_i;
wire na1365_1;
wire na1365_1_i;
wire na1366_1;
wire na1366_1_i;
wire na1367_2;
wire na1367_2_i;
wire na1368_1;
wire na1368_1_i;
wire na1369_1;
wire na1369_1_i;
wire na1370_1;
wire na1370_1_i;
wire na1371_1;
wire na1371_1_i;
wire na1372_1;
wire na1373_1;
wire na1374_2;
wire na1375_2;
wire na1376_2;
wire na1377_1;
wire na1379_1;
wire na1381_1;
wire na1383_1;
wire na1385_1;
wire na1387_1;
wire na1389_1;
wire na1390_2;
wire na1391_2;
wire na1392_1;
wire na1394_1;
wire na1396_1;
wire na1398_1;
wire na1400_1;
wire na1402_1;
wire na1404_1;
wire na1405_1;
wire na1407_1;
wire na1409_1;
wire na1411_1;
wire na1413_1;
wire na1414_1;
wire na1415_1;
wire na1417_1;
wire na1419_1;
wire na1420_2;
wire na1421_1;
wire na1423_1;
wire na1425_1;
wire na1427_1;
wire na1428_1;
wire na1436_1;
wire na1438_1;
wire na1439_1;
wire na1440_1;
wire na1443_1;
wire na1444_1;
wire na1446_1;
wire na1448_1;
wire na1449_1;
wire na1451_1;
wire na1453_1;
wire na1454_1;
wire na1455_1;
wire na1455_1_i;
wire na1456_1;
wire na1457_2;
wire na1458_1;
wire na1459_1;
wire na1460_2;
wire na1461_1;
wire na1462_1;
wire na1464_1;
wire na1465_1;
wire na1466_1;
wire na1467_1;
wire na1469_4;
wire na1471_4;
wire na1473_4;
wire na1474_1;
wire na1474_4;
wire na1475_1;
wire na1475_2;
wire na1475_4;
wire na1477_1;
wire na1477_2;
wire na1477_4;
wire na1479_1;
wire na1479_2;
wire na1481_1;
wire na1481_4;
wire na1482_1;
wire na1482_2;
wire na1482_4;
wire na1484_1;
wire na1487_1;
wire na1487_2;
wire na1488_1;
wire na1488_9;
wire na1489_1;
wire na1489_9;
wire na1592_2;
wire na1592_2_i;
wire na1593_1;
wire na1593_1_i;
wire na1594_2;
wire na1594_2_i;
wire na1595_1;
wire na1595_1_i;
wire na1596_2;
wire na1596_2_i;
wire na1597_1;
wire na1597_1_i;
wire na1598_2;
wire na1598_2_i;
wire na1599_1;
wire na1599_1_i;
wire na1624_2;
wire na1624_2_i;
wire na1625_1;
wire na1625_1_i;
wire na1626_2;
wire na1626_2_i;
wire na1627_1;
wire na1627_1_i;
wire na1628_2;
wire na1628_2_i;
wire na1629_1;
wire na1629_1_i;
wire na1630_2;
wire na1630_2_i;
wire na1631_1;
wire na1631_1_i;
wire na1640_2;
wire na1640_2_i;
wire na1641_1;
wire na1641_1_i;
wire na1642_2;
wire na1642_2_i;
wire na1643_1;
wire na1643_1_i;
wire na1644_2;
wire na1644_2_i;
wire na1645_1;
wire na1645_1_i;
wire na1646_2;
wire na1646_2_i;
wire na1647_1;
wire na1647_1_i;
wire na1648_2;
wire na1648_2_i;
wire na1649_1;
wire na1649_1_i;
wire na1650_2;
wire na1650_2_i;
wire na1651_1;
wire na1651_1_i;
wire na1652_2;
wire na1652_2_i;
wire na1653_1;
wire na1653_1_i;
wire na1654_2;
wire na1654_2_i;
wire na1655_1;
wire na1655_1_i;
wire na1656_2;
wire na1656_2_i;
wire na1657_1;
wire na1657_1_i;
wire na1658_2;
wire na1658_2_i;
wire na1659_1;
wire na1659_1_i;
wire na1660_2;
wire na1660_2_i;
wire na1661_1;
wire na1661_1_i;
wire na1662_2;
wire na1662_2_i;
wire na1663_1;
wire na1663_1_i;
wire na1664_2;
wire na1664_2_i;
wire na1665_1;
wire na1665_1_i;
wire na1666_2;
wire na1666_2_i;
wire na1667_1;
wire na1667_1_i;
wire na1668_2;
wire na1668_2_i;
wire na1669_1;
wire na1669_1_i;
wire na1670_2;
wire na1670_2_i;
wire na1671_1;
wire na1671_1_i;
wire na1672_2;
wire na1672_2_i;
wire na1673_1;
wire na1673_1_i;
wire na1674_2;
wire na1674_2_i;
wire na1675_1;
wire na1675_1_i;
wire na1676_2;
wire na1676_2_i;
wire na1677_1;
wire na1677_1_i;
wire na1678_2;
wire na1678_2_i;
wire na1679_1;
wire na1679_1_i;
wire na1680_2;
wire na1680_2_i;
wire na1681_1;
wire na1681_1_i;
wire na1682_2;
wire na1682_2_i;
wire na1683_1;
wire na1683_1_i;
wire na1684_2;
wire na1684_2_i;
wire na1685_1;
wire na1685_1_i;
wire na1686_2;
wire na1686_2_i;
wire na1687_1;
wire na1687_1_i;
wire na2220_2;
wire na2220_2_i;
wire na2221_1;
wire na2221_1_i;
wire na2222_2;
wire na2222_2_i;
wire na2223_1;
wire na2223_1_i;
wire na2224_2;
wire na2224_2_i;
wire na2225_1;
wire na2225_1_i;
wire na2226_2;
wire na2226_2_i;
wire na2227_1;
wire na2227_1_i;
wire na2228_2;
wire na2228_2_i;
wire na2229_1;
wire na2229_1_i;
wire na2230_2;
wire na2230_2_i;
wire na2231_1;
wire na2231_1_i;
wire na2232_2;
wire na2232_2_i;
wire na2233_1;
wire na2233_1_i;
wire na2234_2;
wire na2234_2_i;
wire na2235_1;
wire na2235_1_i;
wire na2236_2;
wire na2236_2_i;
wire na2237_1;
wire na2237_1_i;
wire na2238_2;
wire na2238_2_i;
wire na2239_1;
wire na2239_1_i;
wire na2240_2;
wire na2240_2_i;
wire na2241_1;
wire na2241_1_i;
wire na2242_2;
wire na2242_2_i;
wire na2243_1;
wire na2243_1_i;
wire na2244_2;
wire na2244_2_i;
wire na2245_1;
wire na2245_1_i;
wire na2246_2;
wire na2246_2_i;
wire na2247_1;
wire na2247_1_i;
wire na2248_2;
wire na2248_2_i;
wire na2249_1;
wire na2249_1_i;
wire na2250_2;
wire na2250_2_i;
wire na2251_1;
wire na2251_1_i;
wire na2348_2;
wire na2348_2_i;
wire na2349_1;
wire na2349_1_i;
wire na2350_2;
wire na2350_2_i;
wire na2351_1;
wire na2351_1_i;
wire na2363_1;
wire na2364_1;
wire na2365_1;
wire na2366_1;
wire na2367_1;
wire na2368_1;
wire na2369_1;
wire na2370_1;
wire na2371_1;
wire na2372_1;
wire na2373_1;
wire na2374_1;
wire na2375_1;
wire na2376_1;
wire na2377_1;
wire na2378_1;
wire na2379_1;
wire na2380_1;
wire na2381_1;
wire na2382_1;
wire na2383_1;
wire na2384_1;
wire na2385_1;
wire na2386_1;
wire na2387_1;
wire na2388_1;
wire na2389_1;
wire na2390_1;
wire na2391_1;
wire na2392_1;
wire na2393_1;
wire na2394_1;
wire na2395_1;
wire na2404_1;
wire na2405_1;
wire na2405_2;
wire na2407_1;
wire na2407_2;
wire na2408_2;
wire na2408_2_i;
wire na2409_1;
wire na2409_2;
wire na2410_1;
wire na2410_2;
wire na2411_1;
wire na2411_4;
wire na2412_1;
wire na2413_1;
wire na2413_2;
wire na2414_1;
wire na2414_2;
wire na2416_2;
wire na2418_1;
wire na2423_1;
wire na2423_2;
wire na2425_2;
wire na2426_1;
wire na2426_2;
wire na2428_1;
wire na2428_2;
wire na2429_1;
wire na2430_1;
wire na2430_2;
wire na2431_1;
wire na2432_1;
wire na2436_2;
wire na2438_1;
wire na2439_1;
wire na2440_1;
wire na2440_2;
wire na2441_1;
wire na2443_2;
wire na2444_2;
wire na2445_1;
wire na2446_1;
wire na2446_2;
wire na2447_1;
wire na2448_1;
wire na2450_2;
wire na2451_1;
wire na2453_1;
wire na2454_2;
wire na2455_1;
wire na2456_2;
wire na2457_1;
wire na2458_1;
wire na2459_1;
wire na2459_2;
wire na2460_2;
wire na2461_1;
wire na2463_1;
wire na2464_1;
wire na2464_2;
wire na2465_1;
wire na2467_1;
wire na2469_1;
wire na2472_1;
wire na2473_1;
wire na2474_1;
wire na2474_2;
wire na2475_2;
wire na2477_1;
wire na2478_2;
wire na2479_1;
wire na2480_1;
wire na2481_2;
wire na2482_1;
wire na2484_2;
wire na2485_1;
wire na2485_2;
wire na2486_1;
wire na2489_1;
wire na2491_1;
wire na2492_1;
wire na2493_2;
wire na2494_1;
wire na2495_1;
wire na2495_2;
wire na2497_1;
wire na2498_2;
wire na2499_1;
wire na2500_1;
wire na2500_2;
wire na2502_1;
wire na2503_1;
wire na2503_2;
wire na2504_1;
wire na2504_2;
wire na2507_1;
wire na2509_2;
wire na2510_1;
wire na2512_1;
wire na2513_2;
wire na2514_1;
wire na2515_1;
wire na2515_2;
wire na2517_1;
wire na2518_1;
wire na2518_2;
wire na2519_2;
wire na2521_1;
wire na2522_1;
wire na2523_2;
wire na2524_1;
wire na2525_1;
wire na2525_2;
wire na2526_1;
wire na2526_2;
wire na2529_1;
wire na2529_2;
wire na2531_1;
wire na2533_2;
wire na2534_1;
wire na2534_2;
wire na2535_1;
wire na2536_1;
wire na2537_1;
wire na2538_1;
wire na2540_2;
wire na2541_1;
wire na2542_1;
wire na2542_2;
wire na2543_1;
wire na2543_2;
wire na2546_1;
wire na2547_1;
wire na2548_2;
wire na2549_1;
wire na2549_2;
wire na2551_1;
wire na2553_1;
wire na2554_1;
wire na2555_1;
wire na2555_2;
wire na2556_1;
wire na2556_2;
wire na2559_1;
wire na2561_2;
wire na2562_1;
wire na2564_1;
wire na2565_1;
wire na2565_2;
wire na2566_1;
wire na2566_2;
wire na2570_1;
wire na2571_1;
wire na2572_1;
wire na2572_2;
wire na2573_1;
wire na2575_1;
wire na2575_2;
wire na2576_1;
wire na2578_1;
wire na2578_2;
wire na2579_1;
wire na2581_1;
wire na2581_2;
wire na2582_1;
wire na2584_1;
wire na2584_2;
wire na2585_1;
wire na2587_1;
wire na2587_2;
wire na2588_1;
wire na2590_1;
wire na2590_2;
wire na2591_1;
wire na2593_1;
wire na2593_2;
wire na2594_1;
wire na2596_1;
wire na2596_2;
wire na2597_1;
wire na2599_1;
wire na2599_2;
wire na2600_1;
wire na2602_1;
wire na2602_2;
wire na2603_1;
wire na2605_1;
wire na2605_2;
wire na2606_1;
wire na2608_1;
wire na2608_2;
wire na2609_1;
wire na2611_1;
wire na2611_2;
wire na2612_1;
wire na2614_1;
wire na2614_2;
wire na2615_1;
wire na2617_1;
wire na2617_2;
wire na2618_1;
wire na2620_1;
wire na2620_2;
wire na2621_1;
wire na2623_1;
wire na2623_2;
wire na2624_1;
wire na2626_1;
wire na2626_2;
wire na2627_1;
wire na2629_1;
wire na2629_2;
wire na2630_1;
wire na2632_1;
wire na2632_2;
wire na2633_1;
wire na2635_1;
wire na2635_2;
wire na2636_1;
wire na2638_1;
wire na2638_2;
wire na2639_1;
wire na2641_1;
wire na2641_2;
wire na2642_1;
wire na2644_1;
wire na2644_2;
wire na2645_1;
wire na2647_1;
wire na2647_2;
wire na2648_1;
wire na2650_1;
wire na2650_2;
wire na2651_1;
wire na2653_1;
wire na2653_2;
wire na2654_1;
wire na2656_1;
wire na2656_2;
wire na2657_1;
wire na2659_1;
wire na2659_2;
wire na2660_1;
wire na2662_1;
wire na2662_2;
wire na2663_1;
wire na2668_2;
wire na2669_1;
wire na2670_2;
wire na2671_1;
wire na2671_2;
wire na2672_1;
wire na2677_2;
wire na2678_2;
wire na2680_1;
wire na2682_2;
wire na2684_1;
wire na2685_1;
wire na2686_2;
wire na2688_1;
wire na2690_2;
wire na2691_1;
wire na2693_1;
wire na2693_2;
wire na2694_1;
wire na2694_2;
wire na2696_2;
wire na2697_1;
wire na2698_2;
wire na2699_1;
wire na2700_2;
wire na2701_1;
wire na2702_2;
wire na2703_1;
wire na2704_2;
wire na2705_1;
wire na2706_1;
wire na2706_2;
wire na2707_2;
wire na2712_2;
wire na2714_1;
wire na2714_2;
wire na2716_1;
wire na2716_2;
wire na2718_1;
wire na2718_2;
wire na2719_2;
wire na2720_1;
wire na2721_2;
wire na2722_1;
wire na2722_2;
wire na2723_1;
wire na2724_1;
wire na2724_2;
wire na2725_2;
wire na2729_1;
wire na2729_2;
wire na2730_1;
wire na2731_2;
wire na2733_1;
wire na2734_2;
wire na2736_1;
wire na2737_2;
wire na2738_1;
wire na2739_2;
wire na2740_1;
wire na2741_2;
wire na2742_1;
wire na2743_2;
wire na2744_1;
wire na2745_2;
wire na2746_1;
wire na2748_1;
wire na2748_2;
wire na2750_1;
wire na2750_2;
wire na2751_1;
wire na2751_2;
wire na2756_2;
wire na2757_1;
wire na2757_2;
wire na2758_1;
wire na2758_2;
wire na2759_1;
wire na2760_2;
wire na2761_1;
wire na2762_2;
wire na2763_1;
wire na2765_2;
wire na2766_1;
wire na2766_2;
wire na2769_1;
wire na2769_2;
wire na2770_1;
wire na2771_2;
wire na2773_1;
wire na2774_2;
wire na2775_1;
wire na2776_2;
wire na2777_1;
wire na2778_2;
wire na2779_1;
wire na2780_2;
wire na2781_1;
wire na2782_2;
wire na2855_1;
wire na2855_2;
wire na2856_1;
wire na2857_2;
wire na2858_1;
wire na2859_2;
wire na2860_1;
wire na2861_2;
wire na2862_1;
wire na2904_2;
wire na2905_1;
wire na2906_1;
wire na2908_2;
wire na2909_1;
wire na2912_1;
wire na2918_2;
wire na2922_1;
wire na2923_1;
wire na2923_2;
wire na2925_1;
wire na2926_2;
wire na2927_1;
wire na2930_1;
wire na2931_2;
wire na2933_1;
wire na2934_1;
wire na2934_2;
wire na2936_2;
wire na2937_1;
wire na2939_2;
wire na2940_1;
wire na2942_1;
wire na2950_2;
wire na2951_1;
wire na2952_2;
wire na2953_2;
wire na2954_2;
wire na2955_2;
wire na2956_2;
wire na2957_2;
wire na2958_2;
wire na2959_2;
wire na2960_2;
wire na2961_2;
wire na2962_2;
wire na2963_2;
wire na2964_2;
wire na2965_2;
wire na2966_2;
wire na2967_2;
wire na2968_2;
wire na2969_2;
wire na2970_2;
wire na2971_2;
wire na2972_2;
wire na2973_2;
wire na2974_2;
wire na2975_2;
wire na2976_2;
wire na2977_2;
wire na2978_2;
wire na2979_2;
wire na2980_2;
wire na2981_2;
wire na2982_2;
wire na2983_2;
wire na2984_2;
wire na2985_2;
wire na2986_2;
wire na2987_2;
wire na2988_2;
wire na2989_2;
wire na2990_2;
wire na2991_2;
wire na2992_2;
wire na2993_2;
wire na2994_2;
wire na2995_2;
wire na2996_2;
wire na2997_2;
wire na2998_2;
wire na2999_2;
wire na3000_2;
wire na3001_2;
wire na3002_2;
wire na3003_2;
wire na3004_2;
wire na3005_2;
wire na3006_2;
wire na3007_2;
wire na3008_2;
wire na3009_2;
wire na3010_2;
wire na3011_2;
wire na3012_2;
wire na3013_2;
wire na3014_2;
wire na3015_2;
wire na3016_2;
wire na3017_2;
wire na3018_2;
wire na3019_2;
wire na3020_2;
wire na3021_2;
wire na3022_2;
wire na3023_2;
wire na3024_2;
wire na3025_2;
wire na3026_2;
wire na3027_2;
wire na3028_2;
wire na3029_2;
wire na3030_2;
wire na3031_2;
wire na3032_2;
wire na3033_2;
wire na3034_2;
wire na3035_2;
wire na3036_2;
wire na3037_2;
wire na3038_2;
wire na3039_2;
wire na3040_2;
wire na3041_2;
wire na3042_2;
wire na3043_2;
wire na3044_2;
wire na3045_2;
wire na3046_2;
wire na3047_2;
wire na3048_2;
wire na3049_2;
wire na3050_2;
wire na3051_2;
wire na3052_2;
wire na3053_2;
wire na3054_2;
wire na3055_2;
wire na3056_2;
wire na3057_2;
wire na3058_2;
wire na3059_2;
wire na3060_2;
wire na3061_2;
wire na3062_2;
wire na3063_2;
wire na3064_2;
wire na3065_2;
wire na3066_2;
wire na3067_2;
wire na3068_2;
wire na3069_2;
wire na3070_2;
wire na3071_2;
wire na3072_2;
wire na3073_2;
wire na3074_2;
wire na3075_2;
wire na3076_2;
wire na3077_2;
wire na3078_2;
wire na3079_2;
wire na3080_2;
wire na3081_2;
wire na3082_2;
wire na3083_2;
wire na3084_2;
wire na3085_2;
wire na3086_2;
wire na3087_2;
wire na3088_2;
wire na3089_2;
wire na3090_2;
wire na3091_2;
wire na3092_2;
wire na3093_2;
wire na3094_2;
wire na3095_2;
wire na3096_2;
wire na3097_2;
wire na3098_2;
wire na3099_2;
wire na3100_2;
wire na3101_2;
wire na3102_2;
wire na3103_2;
wire na3104_2;
wire na3105_2;
wire na3106_2;
wire na3107_2;
wire na3108_2;
wire na3109_2;
wire na3110_2;
wire na3111_2;
wire na3112_2;
wire na3113_2;
wire na3114_2;
wire na3115_2;
wire na3116_2;
wire na3117_2;
wire na3118_2;
wire na3119_2;
wire na3120_2;
wire na3121_2;
wire na3122_2;
wire na3123_2;
wire na3124_2;
wire na3125_2;
wire na3126_2;
wire na3127_2;
wire na3128_2;
wire na3129_2;
wire na3130_2;
wire na3131_2;
wire na3132_2;
wire na3133_2;
wire na3134_2;
wire na3135_2;
wire na3136_2;
wire na3137_2;
wire na3138_2;
wire na3139_2;
wire na3140_2;
wire na3141_2;
wire na3142_2;
wire na3143_2;
wire na3144_2;
wire na3145_2;
wire na3146_2;
wire na3147_2;
wire na3148_2;
wire na3149_2;
wire na3150_2;
wire na3151_2;
wire na3152_2;
wire na3153_2;
wire na3154_2;
wire na3155_2;
wire na3156_2;
wire na3157_2;
wire na3158_2;
wire na3159_2;
wire na3160_2;
wire na3161_2;
wire na3162_2;
wire na3163_2;
wire na3164_2;
wire na3165_2;
wire na3166_2;
wire na3167_2;
wire na3168_2;
wire na3169_2;
wire na3170_2;
wire na3171_2;
wire na3172_2;
wire na3173_2;
wire na3174_2;
wire na3175_2;
wire na3176_2;
wire na3177_2;
wire na3178_2;
wire na3179_2;
wire na3180_2;
wire na3181_2;
wire na3182_2;
wire na3183_2;
wire na3184_2;
wire na3185_2;
wire na3186_2;
wire na3187_2;
wire na3188_2;
wire na3189_2;
wire na3190_2;
wire na3191_2;
wire na3192_2;
wire na3193_2;
wire na3194_2;
wire na3195_2;
wire na3196_2;
wire na3197_2;
wire na3198_2;
wire na3199_2;
wire na3200_2;
wire na3201_2;
wire na3202_2;
wire na3203_2;
wire na3204_2;
wire na3205_2;
wire na3206_2;
wire na3207_2;
wire na3208_2;
wire na3209_2;
wire na3210_2;
wire na3211_2;
wire na3212_2;
wire na3213_2;
wire na3214_2;
wire na3215_2;
wire na3216_2;
wire na3217_2;
wire na3218_2;
wire na3263_1;
wire na3263_2;
wire na3263_3;
wire na3263_6;
wire na2952_10;
wire na2953_10;
wire na2954_10;
wire na2955_10;
wire na2956_10;
wire na2957_10;
wire na2958_10;
wire na2959_10;

// C_AND////      x87y68     80'h00_0018_00_0000_0888_C141
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1), .IN1(~na6_1), .IN2(~na5_1), .IN3(~na8_2), .IN4(na7_1), .IN5(~na6_2), .IN6(~na5_2), .IN7(1'b1), .IN8(na7_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x89y72     80'h00_EE00_80_0000_0C88_F2F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1475_1), .IN6(~na2_1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5_2 ( .OUT(na5_1), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2_i), .IN1(na1479_2), .IN2(~na2_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5_5 ( .OUT(na5_2), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5_2_i) );
// C_AND/D//AND/D      x87y71     80'h00_EE00_80_0000_0C88_F2F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1475_2), .IN6(~na2_1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6_2 ( .OUT(na6_1), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6_4 ( .OUT(na6_2_i), .IN1(na1479_1), .IN2(~na2_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6_5 ( .OUT(na6_2), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_2_i) );
// C_AND/D//AND/D      x88y70     80'h00_EE00_80_0000_0C88_3C33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1477_1), .IN7(1'b1), .IN8(~na2960_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a7_2 ( .OUT(na7_1), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na7_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7_4 ( .OUT(na7_2_i), .IN1(1'b1), .IN2(~na2_1), .IN3(1'b1), .IN4(~na7_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a7_5 ( .OUT(na7_2), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na7_2_i) );
// C_///AND/D      x86y71     80'h00_EE00_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8_4 ( .OUT(na8_2_i), .IN1(1'b1), .IN2(na1477_2), .IN3(1'b1), .IN4(~na2960_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a8_5 ( .OUT(na8_2), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na8_2_i) );
// C_XOR////D      x81y97     80'h40_E818_00_0000_0666_C056
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1), .IN1(~na43_1), .IN2(~na49_1), .IN3(~na37_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na13_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a11_5 ( .OUT(na11_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na11_1) );
// C_ANDXOR////      x80y94     80'h00_0018_00_0000_0666_FE37
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(na2963_2), .IN2(na23_1), .IN3(1'b1), .IN4(na34_1), .IN5(~na2971_2), .IN6(~na23_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y80     80'h00_0018_00_0040_0AF3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1), .IN1(~na1443_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2407_2), .IN5(~na27_1), .IN6(~na2414_2), .IN7(na3173_2),
                    .IN8(na2407_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y105     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3131_2), .IN6(na1031_1), .IN7(na1027_1), .IN8(na1029_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x79y105     80'h00_0018_00_0000_0C88_95FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na20_1), .IN6(1'b0), .IN7(~na1027_1), .IN8(~na3133_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x79y109     80'h00_0078_00_0000_0C66_3AC3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1033_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1021_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a20_4 ( .OUT(na20_2), .IN1(1'b0), .IN2(~na1023_1), .IN3(1'b0), .IN4(na1021_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y108     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2968_2), .IN5(1'b0), .IN6(~na1023_1), .IN7(1'b0), .IN8(~na1021_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x79y98     80'h00_0078_00_0000_0C66_9969
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1033_1), .IN6(na1023_1), .IN7(na1025_1), .IN8(~na1029_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a23_4 ( .OUT(na23_2), .IN1(na1033_1), .IN2(~na1031_1), .IN3(na1027_1), .IN4(na1021_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x82y110     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a25_4 ( .OUT(na25_2), .IN1(~na1033_1), .IN2(na1023_1), .IN3(na1027_1), .IN4(~na1021_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x79y95     80'h00_0018_00_0000_0666_BA57
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(na3168_2), .IN2(na23_1), .IN3(na29_1), .IN4(1'b1), .IN5(~na3132_2), .IN6(1'b1), .IN7(~na2409_2),
                    .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y107     80'h00_0018_00_0040_0AD9_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a29_1 ( .OUT(na29_1), .IN1(1'b1), .IN2(na23_2), .IN3(1'b1), .IN4(~na2410_2), .IN5(~na20_2), .IN6(1'b0), .IN7(na3169_2),
                    .IN8(~na2965_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y104     80'h00_0018_00_0040_0AE1_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1), .IN1(1'b1), .IN2(~na2413_2), .IN3(1'b1), .IN4(~na2410_2), .IN5(1'b1), .IN6(na23_2), .IN7(na1018_1),
                    .IN8(na3172_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y81     80'h00_0018_00_0040_0AF9_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1), .IN1(~na1443_1), .IN2(1'b1), .IN3(~na3173_2), .IN4(1'b1), .IN5(~na27_1), .IN6(na2414_1), .IN7(na2970_2),
                    .IN8(~na2407_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x80y86     80'h00_0018_00_0040_0CA7_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_1 ( .OUT(na34_1), .IN1(na3170_2), .IN2(~na2979_2), .IN3(na2409_2), .IN4(1'b1), .IN5(na2972_2), .IN6(1'b1), .IN7(~na36_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x82y78     80'h00_0018_00_0040_0AF3_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1), .IN1(na27_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2407_2), .IN5(~na1443_1), .IN6(~na3174_2), .IN7(na3173_2),
                    .IN8(na2416_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y81     80'h00_0018_00_0040_0AF8_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(~na27_1), .IN2(1'b1), .IN3(~na3173_2), .IN4(1'b1), .IN5(na1443_1), .IN6(na2418_1), .IN7(na3167_2),
                    .IN8(~na2407_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x82y91     80'h00_0018_00_0000_0666_BF75
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1), .IN1(na38_1), .IN2(1'b1), .IN3(na36_1), .IN4(na2973_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na33_1), .IN8(na2976_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y79     80'h00_0018_00_0040_0AED_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1), .IN1(1'b1), .IN2(na15_1), .IN3(1'b1), .IN4(~na35_1), .IN5(1'b1), .IN6(na2428_2), .IN7(~na1018_1),
                    .IN8(~na45_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x79y73     80'h00_0078_00_0000_0C66_0609
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na20_2), .IN6(na23_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a42_4 ( .OUT(na42_2), .IN1(na20_1), .IN2(~na23_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x79y69     80'h00_0018_00_0000_0666_BF57
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1), .IN1(na42_1), .IN2(na15_1), .IN3(na46_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na33_1), .IN8(na45_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x80y70     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na2428_2), .IN7(na1018_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y71     80'h00_0018_00_0040_0A7E_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1), .IN1(1'b1), .IN2(na3175_2), .IN3(1'b1), .IN4(na35_1), .IN5(na2423_1), .IN6(~na2974_2), .IN7(~na36_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x79y91     80'h00_0078_00_0000_0C66_AC60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1023_1), .IN7(na1025_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a48_4 ( .OUT(na48_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2409_2), .IN4(na2410_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y84     80'h00_0018_00_0000_0666_CC95
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1), .IN1(~na54_1), .IN2(1'b0), .IN3(na50_1), .IN4(~na2426_1), .IN5(1'b0), .IN6(na51_1), .IN7(1'b0), .IN8(na2426_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y89     80'h00_0018_00_0040_0A79_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1), .IN1(1'b1), .IN2(~na15_1), .IN3(1'b1), .IN4(na35_1), .IN5(~na48_2), .IN6(na3171_2), .IN7(na2409_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y86     80'h00_0018_00_0040_0A7E_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1), .IN1(1'b1), .IN2(na23_2), .IN3(na33_1), .IN4(1'b1), .IN5(na2425_2), .IN6(~na23_1), .IN7(~na36_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y95     80'h00_0018_00_0040_0A7C_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1), .IN1(1'b1), .IN2(~na23_1), .IN3(na2969_2), .IN4(1'b1), .IN5(na2972_2), .IN6(na2428_1), .IN7(~na36_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x83y85     80'h40_E800_80_0000_0C88_2F5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2429_1), .IN8(~na2985_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a55_2 ( .OUT(na55_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na55_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a55_4 ( .OUT(na55_2_i), .IN1(1'b1), .IN2(na2479_1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a55_5 ( .OUT(na55_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na55_2_i) );
// C_///OR/      x86y93     80'h00_0060_00_0000_0C0E_FF0B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a57_4 ( .OUT(na57_2), .IN1(na2432_1), .IN2(~na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y100     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1085_1), .IN6(na1084_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x90y96     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1672_2), .IN8(na1592_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x105y84     80'h00_0060_00_0000_0C0E_FF3E
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a62_4 ( .OUT(na62_2), .IN1(na1085_1), .IN2(na1084_1), .IN3(1'b0), .IN4(~na1083_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y88     80'h00_0078_00_0000_0C88_555A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1087_2), .IN6(1'b1), .IN7(~na1103_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a65_4 ( .OUT(na65_2), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x86y87     80'h00_0078_00_0000_0C88_F4F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1087_2), .IN6(na2923_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a66_4 ( .OUT(na66_2), .IN1(~na1085_1), .IN2(~na2436_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x82y106     80'h40_E818_00_0000_0666_9A60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1), .IN1(1'b0), .IN2(1'b0), .IN3(na70_1), .IN4(na2426_2), .IN5(na54_1), .IN6(1'b0), .IN7(~na37_1), .IN8(na2426_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a69_5 ( .OUT(na69_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na69_1) );
// C_XOR////      x78y75     80'h00_0018_00_0000_0666_A669
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1), .IN1(na75_1), .IN2(~na72_1), .IN3(~na1444_1), .IN4(~na2977_2), .IN5(na75_2), .IN6(na51_1), .IN7(na50_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y66     80'h00_0018_00_0000_0666_CA59
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_1 ( .OUT(na72_1), .IN1(na2405_1), .IN2(~na74_1), .IN3(~na73_1), .IN4(1'b0), .IN5(na2405_2), .IN6(1'b0), .IN7(1'b0),
                    .IN8(na34_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x80y65     80'h00_0018_00_0040_0C5E_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1), .IN1(1'b1), .IN2(na2428_1), .IN3(~na36_1), .IN4(na35_1), .IN5(na42_1), .IN6(1'b1), .IN7(na2975_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y64     80'h00_0018_00_0040_0ABC_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1), .IN1(1'b1), .IN2(na15_1), .IN3(na33_1), .IN4(1'b1), .IN5(na2423_2), .IN6(na2438_1), .IN7(1'b1), .IN8(~na45_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x79y67     80'h00_0078_00_0000_0C88_5AF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na42_1), .IN6(1'b1), .IN7(~na33_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a75_4 ( .OUT(na75_2), .IN1(na42_2), .IN2(na15_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x93y83     80'h00_0078_00_0000_0C88_F8F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a82_1 ( .OUT(na82_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1087_2), .IN6(na104_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a82_4 ( .OUT(na82_2), .IN1(~na1087_2), .IN2(na104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y100     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na1593_1), .IN6(na1673_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x83y90     80'h40_E818_00_0000_0666_A0C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1), .IN1(~na88_2), .IN2(1'b0), .IN3(1'b0), .IN4(na86_1), .IN5(1'b0), .IN6(1'b0), .IN7(na70_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a85_5 ( .OUT(na85_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na85_1) );
// C_XOR////      x80y78     80'h00_0018_00_0000_0666_96C6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1), .IN1(na3176_2), .IN2(na49_1), .IN3(1'b0), .IN4(na13_1), .IN5(na54_1), .IN6(na72_1), .IN7(~na37_1),
                    .IN8(na2426_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x77y67     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a88_4 ( .OUT(na88_2), .IN1(~na43_1), .IN2(~na49_1), .IN3(1'b0), .IN4(na13_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x87y87     80'h00_0060_00_0000_0C0E_FFA3
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a91_4 ( .OUT(na91_2), .IN1(1'b0), .IN2(~na104_2), .IN3(na2448_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y88     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na1674_2), .IN6(na1594_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x83y79     80'h40_E818_00_0000_0666_0A60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1), .IN1(1'b0), .IN2(1'b0), .IN3(na95_1), .IN4(na86_1), .IN5(na88_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a94_5 ( .OUT(na94_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na94_1) );
// C_XOR////      x82y69     80'h00_0018_00_0000_0666_096C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a95_1 ( .OUT(na95_1), .IN1(1'b0), .IN2(na74_1), .IN3(na73_1), .IN4(na98_1), .IN5(~na97_1), .IN6(na49_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y71     80'h00_0018_00_0040_0AE5_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1), .IN1(1'b1), .IN2(na15_1), .IN3(~na33_1), .IN4(1'b1), .IN5(1'b1), .IN6(na23_2), .IN7(~na2980_2), .IN8(na2450_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y72     80'h00_0018_00_0040_0AE0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_1 ( .OUT(na98_1), .IN1(~na2972_2), .IN2(1'b1), .IN3(na36_1), .IN4(1'b1), .IN5(1'b0), .IN6(na23_1), .IN7(na2978_2), .IN8(na2451_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x87y80     80'h40_E800_80_0000_0C07_FFB7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a99_4 ( .OUT(na99_2_i), .IN1(~na94_1), .IN2(~na104_1), .IN3(na66_1), .IN4(~na2453_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a99_5 ( .OUT(na99_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na99_2_i) );
// C_MX4b////      x89y83     80'h00_0018_00_0040_0A50_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1), .IN1(1'b1), .IN2(na62_2), .IN3(na3155_2), .IN4(1'b1), .IN5(na1675_1), .IN6(1'b0), .IN7(na1595_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x95y86     80'h00_0078_00_0000_0C88_1F3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na66_2), .IN8(~na2985_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a104_4 ( .OUT(na104_2), .IN1(1'b1), .IN2(na59_1), .IN3(1'b1), .IN4(~na1083_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x87y76     80'h40_E818_00_0000_0666_A0CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1), .IN1(1'b0), .IN2(na106_1), .IN3(1'b0), .IN4(na86_1), .IN5(1'b0), .IN6(1'b0), .IN7(na95_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a105_5 ( .OUT(na105_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na105_1) );
// C_XOR////      x81y70     80'h00_0018_00_0000_0666_06A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1), .IN1(na75_2), .IN2(na72_1), .IN3(na1444_1), .IN4(1'b0), .IN5(na75_1), .IN6(na49_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x82y72     80'h40_E800_80_0000_0C88_5C5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2458_1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a107_2 ( .OUT(na107_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na107_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a107_4 ( .OUT(na107_2_i), .IN1(na2551_1), .IN2(1'b1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a107_5 ( .OUT(na107_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na107_2_i) );
// C_///OR/      x90y79     80'h00_0060_00_0000_0C0E_FFC3
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a109_4 ( .OUT(na109_2), .IN1(1'b0), .IN2(~na104_2), .IN3(1'b0), .IN4(na2461_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x92y78     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na1676_2), .IN6(na1596_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x87y65     80'h40_E818_00_0000_0666_C300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na113_1), .IN7(1'b0), .IN8(na115_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a112_5 ( .OUT(na112_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na112_1) );
// C_XOR////      x81y66     80'h00_0018_00_0000_0666_C6A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1), .IN1(~na43_1), .IN2(na74_1), .IN3(na73_1), .IN4(1'b0), .IN5(~na97_1), .IN6(~na106_1), .IN7(1'b0),
                     .IN8(na98_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x84y64     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a115_1 ( .OUT(na115_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na74_1), .IN7(na73_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x93y71     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na1597_1), .IN6(na1677_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x88y69     80'h00_0060_00_0000_0C0E_FFA3
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a120_4 ( .OUT(na120_2), .IN1(1'b0), .IN2(~na104_2), .IN3(na2467_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x87y67     80'h40_E818_00_0000_0666_0CC0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na122_2), .IN5(1'b0), .IN6(na113_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a121_5 ( .OUT(na121_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na121_1) );
// C_///XOR/      x84y70     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a122_4 ( .OUT(na122_2), .IN1(~na2981_2), .IN2(na72_1), .IN3(na70_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x81y67     80'h40_E800_00_0000_0388_E7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a123_1 ( .OUT(na123_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na121_1), .IN6(~na104_1), .IN7(na66_1), .IN8(na2469_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a123_2 ( .OUT(na123_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na123_1_i) );
// C_MX4b////      x93y75     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na1678_2), .IN6(na1598_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x83y69     80'h40_E818_00_0000_0666_6969
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(na43_1), .IN2(~na106_1), .IN3(na70_1), .IN4(na2990_2), .IN5(~na97_1), .IN6(na74_1), .IN7(na73_1),
                     .IN8(na98_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a128_5 ( .OUT(na128_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na128_1) );
// C_AND/D//AND/D      x82y75     80'h40_E800_80_0000_0C88_5A53
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a129_1 ( .OUT(na129_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2473_1), .IN6(1'b1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a129_2 ( .OUT(na129_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na129_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a129_4 ( .OUT(na129_2_i), .IN1(1'b1), .IN2(~na2546_1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a129_5 ( .OUT(na129_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na129_2_i) );
// C_MX4b////      x91y75     80'h00_0018_00_0040_0AA0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1), .IN1(1'b1), .IN2(~na62_2), .IN3(na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na1679_1), .IN7(1'b0), .IN8(na1599_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y84     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a137_1 ( .OUT(na137_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na977_1), .IN6(na2244_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y82     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na693_2), .IN8(na953_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y87     80'h00_0018_00_0040_0A3F_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a139_1 ( .OUT(na139_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(~na1624_2), .IN6(~na738_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x83y95     80'h40_E800_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na141_1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a140_2 ( .OUT(na140_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na140_1_i) );
// C_AND////      x95y96     80'h00_0018_00_0000_0888_5413
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1), .IN1(1'b1), .IN2(~na144_1), .IN3(~na2485_2), .IN4(~na2482_1), .IN5(~na143_1), .IN6(na2484_2), .IN7(~na2485_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y89     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a143_1 ( .OUT(na143_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na2245_1), .IN6(na978_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y92     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a144_1 ( .OUT(na144_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na954_1), .IN6(na3087_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x82y92     80'h40_E800_80_0000_0C88_5A5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2486_1), .IN6(1'b1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a146_2 ( .OUT(na146_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na146_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a146_4 ( .OUT(na146_2_i), .IN1(1'b1), .IN2(na2439_1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a146_5 ( .OUT(na146_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na146_2_i) );
// C_MX4b////      x98y86     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na2246_2), .IN6(na979_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y87     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a149_1 ( .OUT(na149_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na748_2), .IN6(na955_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y85     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(1'b1), .IN8(na931_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a150_4 ( .OUT(na150_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1666_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y90     80'h00_0018_00_0040_0A3F_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a151_1 ( .OUT(na151_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(~na1626_2), .IN6(~na753_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x82y74     80'h40_E800_80_0000_0C88_2F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2489_1), .IN8(~na2985_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a152_2 ( .OUT(na152_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na152_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a152_4 ( .OUT(na152_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na66_1), .IN4(na2564_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a152_5 ( .OUT(na152_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na152_2_i) );
// C_///AND/      x95y82     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a153_4 ( .OUT(na153_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1667_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y80     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na2247_1), .IN6(na980_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y81     80'h00_0018_00_0040_0A3F_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a156_1 ( .OUT(na156_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(~na1627_1), .IN6(~na759_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y79     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na754_2), .IN6(na956_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y77     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a162_1 ( .OUT(na162_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na66_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2248_2), .IN8(na981_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y76     80'h00_0018_00_0040_0A50_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a163_1 ( .OUT(na163_1), .IN1(1'b1), .IN2(na62_2), .IN3(~na3155_2), .IN4(1'b1), .IN5(na957_1), .IN6(1'b0), .IN7(na760_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x88y65     80'h40_E800_80_0000_0C88_1F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na66_1), .IN8(~na2497_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a164_2 ( .OUT(na164_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na164_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a164_4 ( .OUT(na164_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na66_1), .IN4(na2554_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a164_5 ( .OUT(na164_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na164_2_i) );
// C_MX4b////      x97y70     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na2249_1), .IN6(na982_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y67     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a169_1 ( .OUT(na169_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na958_1), .IN6(na3090_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y72     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na2250_2), .IN6(na983_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y69     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a175_1 ( .OUT(na175_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na769_2), .IN6(na959_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x81y77     80'h40_E800_80_0000_0C88_5C4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a176_1 ( .OUT(na176_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2507_1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a176_2 ( .OUT(na176_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na176_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a176_4 ( .OUT(na176_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na66_1), .IN4(na2445_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a176_5 ( .OUT(na176_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na176_2_i) );
// C_AND///AND/      x97y74     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na936_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a178_4 ( .OUT(na178_2), .IN1(na1631_1), .IN2(1'b1), .IN3(1'b1), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y73     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na66_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2251_1), .IN8(na984_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y71     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na960_1), .IN6(na771_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y96     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na1648_2), .IN6(na985_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y93     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na66_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1649_1), .IN8(na986_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x80y105     80'h40_E800_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a184_4 ( .OUT(na184_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na66_1), .IN4(~na2512_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a184_5 ( .OUT(na184_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na184_2_i) );
// C_MX4b////      x86y104     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na987_1), .IN6(na1650_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x91y105     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a189_1 ( .OUT(na189_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na2238_2), .IN6(na963_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x81y84     80'h40_E800_80_0000_0C88_5A5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a190_1 ( .OUT(na190_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2517_1), .IN6(1'b1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a190_2 ( .OUT(na190_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na190_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a190_4 ( .OUT(na190_2_i), .IN1(1'b1), .IN2(na2541_1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a190_5 ( .OUT(na190_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na190_2_i) );
// C_MX4b////      x87y97     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na1651_1), .IN6(na988_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y97     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2239_1),
                     .IN8(na964_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y100     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a195_4 ( .OUT(na195_2), .IN1(na838_1), .IN2(1'b1), .IN3(1'b1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x85y71     80'h40_E800_80_0000_0C88_4F55
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a196_1 ( .OUT(na196_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na66_1), .IN8(na2521_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a196_2 ( .OUT(na196_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na196_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a196_4 ( .OUT(na196_2_i), .IN1(~na2492_1), .IN2(1'b1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a196_5 ( .OUT(na196_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na196_2_i) );
// C_MX4b////      x91y99     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na1652_2), .IN6(na989_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y100     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a200_1 ( .OUT(na200_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2240_2),
                     .IN8(na965_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y100     80'h00_0018_00_0040_0ACF_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a201_1 ( .OUT(na201_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1660_2),
                     .IN8(~na841_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x83y66     80'h40_E800_80_0000_0C88_2F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2524_1), .IN8(~na2985_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a202_2 ( .OUT(na202_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na202_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a202_4 ( .OUT(na202_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na66_1), .IN4(na2463_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a202_5 ( .OUT(na202_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na202_2_i) );
// C_MX4b////      x112y89     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a205_1 ( .OUT(na205_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na2241_1), .IN6(na966_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y90     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na1653_1), .IN6(na990_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x85y68     80'h40_E800_80_0000_0C88_555A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_1 ( .OUT(na208_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na209_1), .IN6(1'b1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a208_2 ( .OUT(na208_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na208_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a208_4 ( .OUT(na208_2_i), .IN1(na2502_1), .IN2(1'b1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a208_5 ( .OUT(na208_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na208_2_i) );
// C_AND////      x103y85     80'h00_0018_00_0000_0888_43F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a209_1 ( .OUT(na209_1), .IN1(~na3180_2), .IN2(~na211_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2529_1), .IN7(~na212_1),
                     .IN8(na213_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y86     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a211_1 ( .OUT(na211_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na2242_2), .IN6(na967_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y87     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na1654_2), .IN6(na991_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y88     80'h00_0018_00_0040_0A3F_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a213_1 ( .OUT(na213_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(~na1662_2), .IN6(~na846_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x82y81     80'h40_E800_80_0000_0C88_555A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na215_1), .IN6(1'b1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a214_2 ( .OUT(na214_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na214_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a214_4 ( .OUT(na214_2_i), .IN1(na1449_1), .IN2(1'b1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a214_5 ( .OUT(na214_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na214_2_i) );
// C_AND////      x95y99     80'h00_0018_00_0000_0888_1A31
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a215_1 ( .OUT(na215_1), .IN1(~na2531_1), .IN2(~na217_1), .IN3(1'b1), .IN4(~na2534_2), .IN5(na2533_2), .IN6(1'b1), .IN7(~na218_1),
                     .IN8(~na2534_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y96     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a217_1 ( .OUT(na217_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na66_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1655_1), .IN8(na992_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y97     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na2243_1), .IN6(na968_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x84y90     80'h40_E800_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na66_1), .IN8(na2535_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a220_2 ( .OUT(na220_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na220_1_i) );
// C_MX4b////      x89y96     80'h00_0018_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a223_1 ( .OUT(na223_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(~na66_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na993_1), .IN8(na1680_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x94y96     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na969_1), .IN6(na1640_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x88y97     80'h00_0018_00_0040_0A3F_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_1 ( .OUT(na225_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(~na849_2), .IN6(~na898_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x83y95     80'h40_E800_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a226_4 ( .OUT(na226_2_i), .IN1(na2538_1), .IN2(1'b1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a226_5 ( .OUT(na226_2), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na226_2_i) );
// C_///AND/      x90y107     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a227_4 ( .OUT(na227_2), .IN1(na82_2), .IN2(na2229_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y102     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na994_1), .IN6(na1681_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y107     80'h00_0018_00_0040_0ACF_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a230_1 ( .OUT(na230_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na907_1),
                     .IN8(~na899_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y105     80'h00_0018_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na970_1),
                     .IN8(na1641_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y100     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_1 ( .OUT(na235_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na1642_2), .IN6(na971_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x88y99     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na995_1), .IN6(na1682_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x90y91     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a242_1 ( .OUT(na242_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na1683_1), .IN6(na996_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y90     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na972_1), .IN6(na1643_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y87     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a245_1 ( .OUT(na245_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2232_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x91y86     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_1 ( .OUT(na247_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na997_1), .IN6(na1684_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y91     80'h00_0018_00_0040_0ACF_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a248_1 ( .OUT(na248_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na918_2),
                     .IN8(~na920_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y87     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1644_2),
                     .IN8(na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y81     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a253_1 ( .OUT(na253_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na998_1), .IN6(na1685_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y81     80'h00_0018_00_0040_0AA0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a255_1 ( .OUT(na255_1), .IN1(1'b1), .IN2(~na62_2), .IN3(~na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na974_1), .IN7(1'b0), .IN8(na1645_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x82y66     80'h40_E800_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2559_1), .IN6(1'b1), .IN7(~na66_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a256_2 ( .OUT(na256_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na256_1_i) );
// C_AND///AND/      x95y74     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_1 ( .OUT(na258_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na951_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a258_4 ( .OUT(na258_2), .IN1(na925_2), .IN2(1'b1), .IN3(1'b1), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y75     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na66_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1686_2), .IN8(na999_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y75     80'h00_0018_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a261_1 ( .OUT(na261_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na975_1),
                     .IN8(na1646_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x93y82     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na66_2), .IN4(1'b1), .IN5(na1687_1), .IN6(na1000_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y81     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na976_1), .IN6(na1647_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x92y98     80'h40_E800_00_0000_0788_3B57
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a268_1 ( .OUT(na268_1_i), .IN1(~na2570_1), .IN2(~na104_1), .IN3(~na272_1), .IN4(1'b0), .IN5(na2571_1), .IN6(~na104_2), .IN7(1'b0),
                     .IN8(~na271_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a268_2 ( .OUT(na268_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na268_1_i) );
// C_MX4b////      x94y100     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_1 ( .OUT(na271_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na3010_2), .IN6(na469_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x92y101     80'h00_0018_00_0040_0AA0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1), .IN1(1'b1), .IN2(~na62_2), .IN3(~na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na3053_2), .IN7(1'b0), .IN8(na525_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x82y105     80'h40_E800_00_0000_0EEE_E0CE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1_i), .IN1(na277_1), .IN2(na276_1), .IN3(1'b0), .IN4(na2572_2), .IN5(1'b0), .IN6(1'b0), .IN7(na274_1),
                     .IN8(na2572_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a273_2 ( .OUT(na273_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na273_1_i) );
// C_AND////      x86y99     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a274_1 ( .OUT(na274_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na104_1), .IN7(1'b1), .IN8(na2573_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y104     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na430_1), .IN6(na470_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y103     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na526_2), .IN8(na3054_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x86y95     80'h40_E800_00_0000_0EEE_E0CE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1_i), .IN1(na281_1), .IN2(na282_1), .IN3(1'b0), .IN4(na2575_2), .IN5(1'b0), .IN6(1'b0), .IN7(na279_2),
                     .IN8(na2575_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a278_2 ( .OUT(na278_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na278_1_i) );
// C_///AND/      x88y91     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a279_4 ( .OUT(na279_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2576_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x91y91     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a281_1 ( .OUT(na281_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3014_2),
                     .IN8(na471_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x89y94     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na623_1), .IN6(na527_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x88y81     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1_i), .IN1(na286_1), .IN2(na287_1), .IN3(na2578_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2578_1),
                     .IN8(na284_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a283_2 ( .OUT(na283_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na283_1_i) );
// C_AND////      x90y82     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2579_1), .IN6(na104_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x91y81     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a286_1 ( .OUT(na286_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na432_2), .IN6(na3031_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x93y80     80'h00_0018_00_0040_0AA0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1), .IN1(1'b1), .IN2(~na62_2), .IN3(~na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na3055_2), .IN7(1'b0), .IN8(na528_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y68     80'h40_E800_00_0000_0EEE_CCEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_1 ( .OUT(na288_1_i), .IN1(1'b0), .IN2(na292_1), .IN3(na291_1), .IN4(na2581_2), .IN5(1'b0), .IN6(na289_2), .IN7(1'b0),
                     .IN8(na2581_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a288_2 ( .OUT(na288_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na288_1_i) );
// C_///AND/      x91y72     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a289_4 ( .OUT(na289_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2582_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x94y75     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a291_1 ( .OUT(na291_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na473_2), .IN6(na3015_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y70     80'h00_0018_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a292_1 ( .OUT(na292_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na3056_2),
                     .IN8(na529_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x98y66     80'h40_E800_00_0000_0EEE_CACE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a293_1 ( .OUT(na293_1_i), .IN1(na297_1), .IN2(na296_1), .IN3(1'b0), .IN4(na2584_2), .IN5(na294_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na2584_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a293_2 ( .OUT(na293_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na293_1_i) );
// C_///AND/      x95y69     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a294_4 ( .OUT(na294_2), .IN1(1'b1), .IN2(na104_1), .IN3(na2585_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y70     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a296_1 ( .OUT(na296_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3016_2),
                     .IN8(na474_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y67     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a297_1 ( .OUT(na297_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na530_1), .IN6(na3057_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x95y67     80'h40_E800_00_0000_0EEE_CECA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a298_1 ( .OUT(na298_1_i), .IN1(na301_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2587_2), .IN5(na302_1), .IN6(na299_2), .IN7(1'b0),
                     .IN8(na2587_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a298_2 ( .OUT(na298_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na298_1_i) );
// C_///AND/      x91y70     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a299_4 ( .OUT(na299_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2588_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y71     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a301_1 ( .OUT(na301_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na435_1), .IN6(na3033_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x97y67     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a302_1 ( .OUT(na302_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na531_1), .IN8(na627_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x96y67     80'h40_E800_00_0000_0EEE_ACEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a303_1 ( .OUT(na303_1_i), .IN1(1'b0), .IN2(na2590_2), .IN3(na307_1), .IN4(na306_1), .IN5(1'b0), .IN6(na2590_1), .IN7(na304_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a303_2 ( .OUT(na303_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na303_1_i) );
// C_///AND/      x94y71     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a304_4 ( .OUT(na304_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2591_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y74     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a306_1 ( .OUT(na306_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na436_2), .IN6(na476_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y69     80'h00_0018_00_0040_0AA0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_1 ( .OUT(na307_1), .IN1(1'b1), .IN2(~na62_2), .IN3(~na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na628_1), .IN7(1'b0), .IN8(na532_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x112y94     80'h40_E800_00_0000_0EEE_AAAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a308_1 ( .OUT(na308_1_i), .IN1(na2593_2), .IN2(na312_1), .IN3(na311_1), .IN4(1'b0), .IN5(na2593_1), .IN6(1'b0), .IN7(na309_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a308_2 ( .OUT(na308_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na308_1_i) );
// C_AND////      x106y89     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na104_1), .IN7(na2594_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y93     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na437_2), .IN6(na477_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y96     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_1 ( .OUT(na312_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na629_2), .IN6(na533_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x103y105     80'h40_E800_00_0000_0EEE_CCEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a313_1 ( .OUT(na313_1_i), .IN1(na317_1), .IN2(1'b0), .IN3(na316_1), .IN4(na2596_2), .IN5(1'b0), .IN6(na314_2), .IN7(1'b0),
                     .IN8(na2596_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a313_2 ( .OUT(na313_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na313_1_i) );
// C_///AND/      x105y98     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a314_4 ( .OUT(na314_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2597_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y105     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_1 ( .OUT(na316_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na438_1), .IN8(na478_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y103     80'h00_0018_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a317_1 ( .OUT(na317_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na630_1),
                     .IN8(na534_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x116y86     80'h40_E800_00_0000_0EEE_E0EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_1 ( .OUT(na318_1_i), .IN1(na322_1), .IN2(1'b0), .IN3(na321_1), .IN4(na2599_2), .IN5(1'b0), .IN6(1'b0), .IN7(na319_1),
                     .IN8(na2599_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a318_2 ( .OUT(na318_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na318_1_i) );
// C_AND////      x112y85     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2600_1), .IN6(na104_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y87     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na439_2), .IN8(na3038_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y83     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na535_1), .IN6(na3058_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x112y79     80'h40_E800_00_0000_0EEE_CCCE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a323_1 ( .OUT(na323_1_i), .IN1(na327_1), .IN2(na326_1), .IN3(1'b0), .IN4(na2602_2), .IN5(1'b0), .IN6(na324_1), .IN7(1'b0),
                     .IN8(na2602_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a323_2 ( .OUT(na323_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na323_1_i) );
// C_AND////      x107y78     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na104_1), .IN7(na2603_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y82     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a326_1 ( .OUT(na326_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na440_1), .IN6(na480_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y79     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na536_2), .IN8(na632_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x109y73     80'h40_E800_00_0000_0EEE_E0EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1_i), .IN1(na332_1), .IN2(1'b0), .IN3(na2605_2), .IN4(na331_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2605_1),
                     .IN8(na329_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a328_2 ( .OUT(na328_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na328_1_i) );
// C_AND////      x106y78     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na104_1), .IN7(1'b1), .IN8(na2606_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y80     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a331_1 ( .OUT(na331_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na481_2), .IN6(na3018_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y77     80'h00_0018_00_0040_0A50_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a332_1 ( .OUT(na332_1), .IN1(1'b1), .IN2(na62_2), .IN3(na3155_2), .IN4(1'b1), .IN5(na537_1), .IN6(1'b0), .IN7(na633_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x110y67     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a333_1 ( .OUT(na333_1_i), .IN1(na336_1), .IN2(na337_1), .IN3(na2608_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2608_1),
                     .IN8(na334_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a333_2 ( .OUT(na333_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na333_1_i) );
// C_///AND/      x102y70     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a334_4 ( .OUT(na334_2), .IN1(1'b1), .IN2(na104_1), .IN3(na2609_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y73     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a336_1 ( .OUT(na336_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na442_1), .IN8(na482_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y74     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a337_1 ( .OUT(na337_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na538_2), .IN8(na634_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x107y70     80'h40_E800_00_0000_0EEE_0EAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a338_1 ( .OUT(na338_1_i), .IN1(na2611_2), .IN2(na341_1), .IN3(na342_1), .IN4(1'b0), .IN5(na2611_1), .IN6(na339_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a338_2 ( .OUT(na338_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na338_1_i) );
// C_///AND/      x103y76     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a339_4 ( .OUT(na339_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2612_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y76     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a341_1 ( .OUT(na341_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na483_2), .IN6(na443_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y71     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a342_1 ( .OUT(na342_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na539_2), .IN6(na635_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x114y70     80'h40_E800_00_0000_0EEE_CAEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1_i), .IN1(na347_1), .IN2(1'b0), .IN3(na346_1), .IN4(na2614_2), .IN5(na344_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na2614_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a343_2 ( .OUT(na343_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na343_1_i) );
// C_///AND/      x105y77     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a344_4 ( .OUT(na344_2), .IN1(1'b1), .IN2(na2615_1), .IN3(1'b1), .IN4(na2992_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y75     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a346_1 ( .OUT(na346_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na444_2), .IN6(na484_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y73     80'h00_0018_00_0040_0AA0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_1 ( .OUT(na347_1), .IN1(1'b1), .IN2(~na62_2), .IN3(na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na540_1), .IN7(1'b0), .IN8(na636_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x114y83     80'h40_E800_00_0000_0EEE_ACAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_1 ( .OUT(na348_1_i), .IN1(na351_1), .IN2(na2617_2), .IN3(na352_1), .IN4(1'b0), .IN5(1'b0), .IN6(na2617_1), .IN7(na349_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a348_2 ( .OUT(na348_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na348_1_i) );
// C_AND////      x112y83     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2618_1), .IN6(na104_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y85     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na3020_2), .IN6(na485_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y81     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na3046_2),
                     .IN8(na637_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x110y79     80'h40_E800_00_0000_0EEE_CCEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1_i), .IN1(1'b0), .IN2(na356_1), .IN3(na357_1), .IN4(na2620_2), .IN5(1'b0), .IN6(na354_1), .IN7(1'b0),
                     .IN8(na2620_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a353_2 ( .OUT(na353_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na353_1_i) );
// C_AND////      x105y80     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na104_1), .IN7(na2621_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y86     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na446_2), .IN6(na486_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y77     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na542_2), .IN8(na638_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x98y109     80'h40_E800_00_0000_0EEE_ACAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a358_1 ( .OUT(na358_1_i), .IN1(na362_1), .IN2(na361_1), .IN3(na2623_2), .IN4(1'b0), .IN5(1'b0), .IN6(na359_1), .IN7(na2623_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a358_2 ( .OUT(na358_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na358_1_i) );
// C_AND////      x97y104     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na104_1), .IN7(1'b1), .IN8(na2624_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y106     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a361_1 ( .OUT(na361_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na447_1), .IN6(na487_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y103     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na639_2), .IN6(na543_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x108y98     80'h40_E800_00_0000_0EEE_CAEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1_i), .IN1(1'b0), .IN2(na366_1), .IN3(na367_1), .IN4(na2626_2), .IN5(na364_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na2626_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a363_2 ( .OUT(na363_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na363_1_i) );
// C_///AND/      x105y95     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a364_4 ( .OUT(na364_2), .IN1(na2627_1), .IN2(na104_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y94     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3021_2),
                     .IN8(na488_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x112y97     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_1 ( .OUT(na367_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na640_1), .IN6(na3047_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x100y107     80'h40_E800_00_0000_0EEE_EAAC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_1 ( .OUT(na368_1_i), .IN1(1'b0), .IN2(na371_1), .IN3(na372_1), .IN4(1'b0), .IN5(na3183_2), .IN6(1'b0), .IN7(na2629_1),
                     .IN8(na369_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a368_2 ( .OUT(na368_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na368_1_i) );
// C_///AND/      x100y98     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a369_4 ( .OUT(na369_2), .IN1(1'b1), .IN2(na104_1), .IN3(na2630_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x101y102     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a371_1 ( .OUT(na371_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na3041_2), .IN6(na449_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y101     80'h00_0018_00_0040_0A50_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a372_1 ( .OUT(na372_1), .IN1(1'b1), .IN2(na62_2), .IN3(na3155_2), .IN4(1'b1), .IN5(na545_1), .IN6(1'b0), .IN7(na641_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x115y88     80'h40_E800_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a373_1 ( .OUT(na373_1_i), .IN1(1'b0), .IN2(na377_1), .IN3(na376_1), .IN4(na2632_2), .IN5(1'b0), .IN6(1'b0), .IN7(na374_2),
                     .IN8(na2632_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a373_2 ( .OUT(na373_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na373_1_i) );
// C_///AND/      x110y85     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a374_4 ( .OUT(na374_2), .IN1(na2633_1), .IN2(na104_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y89     80'h00_0018_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a376_1 ( .OUT(na376_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na490_1),
                     .IN8(na3022_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y88     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a377_1 ( .OUT(na377_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na3048_2),
                     .IN8(na642_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x113y76     80'h40_E800_00_0000_0EEE_ACEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1_i), .IN1(na382_1), .IN2(1'b0), .IN3(na2635_2), .IN4(na381_1), .IN5(1'b0), .IN6(na379_1), .IN7(na2635_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a378_2 ( .OUT(na378_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na378_1_i) );
// C_AND////      x109y76     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_1 ( .OUT(na379_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2636_1), .IN7(1'b1), .IN8(na2992_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x110y78     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na491_2), .IN6(na451_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y75     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_1 ( .OUT(na382_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na547_1), .IN8(na643_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x104y104     80'h40_E800_00_0000_0EEE_AAEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a383_1 ( .OUT(na383_1_i), .IN1(na2638_2), .IN2(1'b0), .IN3(na386_1), .IN4(na387_1), .IN5(na2638_1), .IN6(1'b0), .IN7(na384_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a383_2 ( .OUT(na383_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na383_1_i) );
// C_///AND/      x104y95     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a384_4 ( .OUT(na384_2), .IN1(na2639_1), .IN2(na104_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y99     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na452_1), .IN8(na492_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x108y100     80'h00_0018_00_0040_0AA0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a387_1 ( .OUT(na387_1), .IN1(1'b1), .IN2(~na62_2), .IN3(na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na548_2), .IN7(1'b0), .IN8(na3059_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x94y93     80'h40_E800_00_0000_0EEE_E0CE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a388_1 ( .OUT(na388_1_i), .IN1(na392_1), .IN2(na391_1), .IN3(1'b0), .IN4(na2641_2), .IN5(1'b0), .IN6(1'b0), .IN7(na389_1),
                     .IN8(na2641_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a388_2 ( .OUT(na388_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na388_1_i) );
// C_AND////      x92y89     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a389_1 ( .OUT(na389_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2642_1), .IN6(na104_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y94     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na453_1), .IN8(na461_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y89     80'h00_0018_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a392_1 ( .OUT(na392_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na645_2),
                     .IN8(na549_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x88y107     80'h40_E800_00_0000_0EEE_CAEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1_i), .IN1(1'b0), .IN2(na396_1), .IN3(na397_1), .IN4(na2644_2), .IN5(na394_1), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na2644_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a393_2 ( .OUT(na393_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na393_1_i) );
// C_AND////      x93y103     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a394_1 ( .OUT(na394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2645_1), .IN7(1'b1), .IN8(na2992_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x95y106     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_1 ( .OUT(na396_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na454_2), .IN6(na462_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y105     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a397_1 ( .OUT(na397_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na646_1), .IN6(na550_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y104     80'h40_E800_00_0000_0EEE_CCEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a398_1 ( .OUT(na398_1_i), .IN1(na401_1), .IN2(1'b0), .IN3(na402_1), .IN4(na2647_2), .IN5(1'b0), .IN6(na399_1), .IN7(1'b0),
                     .IN8(na2647_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a398_2 ( .OUT(na398_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na398_1_i) );
// C_AND////      x95y98     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2648_1), .IN7(1'b1), .IN8(na2992_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x93y101     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a401_1 ( .OUT(na401_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na463_2), .IN6(na3026_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x94y101     80'h00_0018_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a402_1 ( .OUT(na402_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na647_2),
                     .IN8(na551_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x102y93     80'h40_E800_00_0000_0EEE_CAAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1_i), .IN1(na2650_1), .IN2(na407_1), .IN3(na406_1), .IN4(1'b0), .IN5(na2650_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na404_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a403_2 ( .OUT(na403_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na403_1_i) );
// C_///AND/      x100y90     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a404_4 ( .OUT(na404_2), .IN1(na2651_1), .IN2(na104_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x102y91     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a406_1 ( .OUT(na406_1), .IN1(na1087_2), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na456_2), .IN8(na3030_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y90     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a407_1 ( .OUT(na407_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na648_1), .IN6(na552_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x106y85     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1_i), .IN1(na411_1), .IN2(na412_1), .IN3(na2653_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2653_1),
                     .IN8(na409_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a408_2 ( .OUT(na408_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na408_1_i) );
// C_///AND/      x102y86     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a409_4 ( .OUT(na409_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2654_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x107y87     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na457_1), .IN6(na465_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y84     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a412_1 ( .OUT(na412_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2982_2), .IN5(1'b0), .IN6(1'b0), .IN7(na553_1), .IN8(na649_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x109y68     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1_i), .IN1(na417_1), .IN2(na416_1), .IN3(na2656_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2656_1),
                     .IN8(na414_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a413_2 ( .OUT(na413_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na413_1_i) );
// C_///AND/      x104y76     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a414_4 ( .OUT(na414_2), .IN1(1'b1), .IN2(na104_1), .IN3(1'b1), .IN4(na2657_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y76     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na466_1), .IN6(na3027_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y69     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na554_2), .IN6(na650_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x100y66     80'h40_E800_00_0000_0EEE_ECAC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a418_1 ( .OUT(na418_1_i), .IN1(1'b0), .IN2(na2659_2), .IN3(na421_1), .IN4(1'b0), .IN5(1'b0), .IN6(na2659_1), .IN7(na422_1),
                     .IN8(na419_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a418_2 ( .OUT(na418_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na418_1_i) );
// C_AND////      x100y72     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a419_1 ( .OUT(na419_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2660_1), .IN7(1'b1), .IN8(na2992_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y73     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na459_2), .IN6(na467_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x104y69     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a422_1 ( .OUT(na422_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(na651_2), .IN6(na555_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x105y71     80'h40_E800_00_0000_0EEE_E0AE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1_i), .IN1(na427_1), .IN2(na426_1), .IN3(na2662_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2662_1),
                     .IN8(na424_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a423_2 ( .OUT(na423_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na423_1_i) );
// C_AND////      x102y76     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a424_1 ( .OUT(na424_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2663_1), .IN7(1'b1), .IN8(na2992_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x109y80     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a426_1 ( .OUT(na426_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(na460_2), .IN6(na468_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y73     80'h00_0018_00_0040_0AA0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_1 ( .OUT(na427_1), .IN1(1'b1), .IN2(~na62_2), .IN3(na3155_2), .IN4(1'b1), .IN5(1'b0), .IN6(na556_2), .IN7(1'b0), .IN8(na652_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x88y101     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a428_1 ( .OUT(na428_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1212_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a428_2 ( .OUT(na428_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na428_1_i) );
// C_OR////      x104y86     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1085_1), .IN6(~na2436_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x83y107     80'h40_E800_80_0000_0C88_4F3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_1 ( .OUT(na430_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1213_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a430_2 ( .OUT(na430_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na430_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a430_4 ( .OUT(na430_2_i), .IN1(1'b1), .IN2(na1125_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a430_5 ( .OUT(na430_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na430_2_i) );
// C_AND/D///      x85y94     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1214_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a431_2 ( .OUT(na431_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na431_1_i) );
// C_///AND/D      x91y87     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a432_4 ( .OUT(na432_2_i), .IN1(1'b1), .IN2(na1215_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a432_5 ( .OUT(na432_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na432_2_i) );
// C_AND/D///      x91y71     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a433_1 ( .OUT(na433_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1216_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a433_2 ( .OUT(na433_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na433_1_i) );
// C_///AND/D      x101y72     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a434_4 ( .OUT(na434_2_i), .IN1(na1217_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a434_5 ( .OUT(na434_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na434_2_i) );
// C_AND/D///      x95y69     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1218_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a435_2 ( .OUT(na435_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na435_1_i) );
// C_///AND/D      x93y69     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a436_4 ( .OUT(na436_2_i), .IN1(na1219_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a436_5 ( .OUT(na436_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na436_2_i) );
// C_///AND/D      x113y93     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a437_4 ( .OUT(na437_2_i), .IN1(na1220_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a437_5 ( .OUT(na437_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na437_2_i) );
// C_AND/D//AND/D      x106y107     80'h40_E800_80_0000_0C88_4F3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1221_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a438_2 ( .OUT(na438_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na438_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a438_4 ( .OUT(na438_2_i), .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a438_5 ( .OUT(na438_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na438_2_i) );
// C_///AND/D      x118y85     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a439_4 ( .OUT(na439_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1222_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a439_5 ( .OUT(na439_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na439_2_i) );
// C_AND/D///      x113y79     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_1 ( .OUT(na440_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1223_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a440_2 ( .OUT(na440_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na440_1_i) );
// C_///AND/D      x114y74     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a441_4 ( .OUT(na441_2_i), .IN1(na1224_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a441_5 ( .OUT(na441_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na441_2_i) );
// C_AND/D///      x112y69     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1225_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a442_2 ( .OUT(na442_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na442_1_i) );
// C_///AND/D      x109y70     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a443_4 ( .OUT(na443_2_i), .IN1(1'b1), .IN2(na1226_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a443_5 ( .OUT(na443_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na443_2_i) );
// C_///AND/D      x113y69     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a444_4 ( .OUT(na444_2_i), .IN1(na1227_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a444_5 ( .OUT(na444_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na444_2_i) );
// C_AND/D///      x120y86     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a445_1 ( .OUT(na445_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1228_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a445_2 ( .OUT(na445_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na445_1_i) );
// C_///AND/D      x117y87     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a446_4 ( .OUT(na446_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1229_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a446_5 ( .OUT(na446_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na446_2_i) );
// C_AND/D///      x105y105     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a447_1 ( .OUT(na447_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1230_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a447_2 ( .OUT(na447_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na447_1_i) );
// C_///AND/D      x115y93     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a448_4 ( .OUT(na448_2_i), .IN1(1'b1), .IN2(na1231_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a448_5 ( .OUT(na448_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na448_2_i) );
// C_AND/D///      x107y104     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_1 ( .OUT(na449_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1232_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a449_2 ( .OUT(na449_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na449_1_i) );
// C_AND/D//AND/D      x118y89     80'h40_E800_80_0000_0C88_4F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a450_1 ( .OUT(na450_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1233_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a450_2 ( .OUT(na450_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na450_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3011_2), .IN4(na1145_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a450_5 ( .OUT(na450_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na450_2_i) );
// C_AND/D///      x115y76     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1234_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a451_2 ( .OUT(na451_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na451_1_i) );
// C_AND/D//AND/D      x110y105     80'h40_E800_80_0000_0C88_4F3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1235_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a452_2 ( .OUT(na452_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na452_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a452_4 ( .OUT(na452_2_i), .IN1(1'b1), .IN2(na1147_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a452_5 ( .OUT(na452_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na452_2_i) );
// C_AND/D///      x102y89     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a453_1 ( .OUT(na453_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1236_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a453_2 ( .OUT(na453_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na453_1_i) );
// C_///AND/D      x99y105     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a454_4 ( .OUT(na454_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1237_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a454_5 ( .OUT(na454_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na454_2_i) );
// C_AND/D///      x100y103     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1238_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a455_2 ( .OUT(na455_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na455_1_i) );
// C_///AND/D      x108y91     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a456_4 ( .OUT(na456_2_i), .IN1(1'b1), .IN2(na1239_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a456_5 ( .OUT(na456_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na456_2_i) );
// C_AND/D///      x115y87     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_1 ( .OUT(na457_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1240_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a457_2 ( .OUT(na457_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na457_1_i) );
// C_///AND/D      x116y76     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a458_4 ( .OUT(na458_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1241_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a458_5 ( .OUT(na458_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na458_2_i) );
// C_///AND/D      x101y73     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a459_4 ( .OUT(na459_2_i), .IN1(1'b1), .IN2(na1242_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a459_5 ( .OUT(na459_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na459_2_i) );
// C_///AND/D      x109y83     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a460_4 ( .OUT(na460_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1243_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a460_5 ( .OUT(na460_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na460_2_i) );
// C_AND/D//AND/D      x86y98     80'h40_E800_80_0000_0C88_3C2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_1 ( .OUT(na461_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1364_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a461_2 ( .OUT(na461_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na461_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a461_4 ( .OUT(na461_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1268_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a461_5 ( .OUT(na461_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na461_2_i) );
// C_AND/D//AND/D      x93y108     80'h40_E800_80_0000_0C88_4F3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a462_1 ( .OUT(na462_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1365_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a462_2 ( .OUT(na462_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na462_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a462_4 ( .OUT(na462_2_i), .IN1(1'b1), .IN2(na1269_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a462_5 ( .OUT(na462_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na462_2_i) );
// C_///AND/D      x93y103     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a463_4 ( .OUT(na463_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1366_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a463_5 ( .OUT(na463_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na463_2_i) );
// C_///AND/D      x103y92     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a464_4 ( .OUT(na464_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1367_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a464_5 ( .OUT(na464_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na464_2_i) );
// C_AND/D///      x107y84     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1368_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a465_2 ( .OUT(na465_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na465_1_i) );
// C_AND/D///      x109y71     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1369_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a466_2 ( .OUT(na466_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na466_1_i) );
// C_AND/D//AND/D      x101y68     80'h40_E800_80_0000_0C88_3C4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1370_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a467_2 ( .OUT(na467_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na467_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a467_4 ( .OUT(na467_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3011_2), .IN4(na1274_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a467_5 ( .OUT(na467_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na467_2_i) );
// C_AND/D//AND/D      x105y70     80'h40_E800_80_0000_0C88_3A4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a468_1 ( .OUT(na468_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1371_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a468_2 ( .OUT(na468_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na468_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a468_4 ( .OUT(na468_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3011_2), .IN4(na1275_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a468_5 ( .OUT(na468_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na468_2_i) );
// C_///AND/D      x93y102     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a469_4 ( .OUT(na469_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1340_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a469_5 ( .OUT(na469_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na469_2_i) );
// C_AND/D//AND/D      x85y106     80'h40_E800_80_0000_0C88_3A3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a470_2 ( .OUT(na470_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na470_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a470_4 ( .OUT(na470_2_i), .IN1(na1245_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a470_5 ( .OUT(na470_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na470_2_i) );
// C_AND/D///      x92y86     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_1 ( .OUT(na471_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1342_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a471_2 ( .OUT(na471_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na471_1_i) );
// C_///AND/D      x92y86     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a472_4 ( .OUT(na472_2_i), .IN1(1'b1), .IN2(na1343_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a472_5 ( .OUT(na472_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na472_2_i) );
// C_///AND/D      x91y69     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a473_4 ( .OUT(na473_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1344_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a473_5 ( .OUT(na473_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na473_2_i) );
// C_///AND/D      x102y68     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a474_4 ( .OUT(na474_2_i), .IN1(na1345_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a474_5 ( .OUT(na474_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na474_2_i) );
// C_AND/D///      x93y65     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_1 ( .OUT(na475_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1346_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a475_2 ( .OUT(na475_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na475_1_i) );
// C_AND/D///      x99y68     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_1 ( .OUT(na476_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1347_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a476_2 ( .OUT(na476_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na476_1_i) );
// C_AND/D///      x119y94     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1348_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a477_2 ( .OUT(na477_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na477_1_i) );
// C_AND/D//AND/D      x108y104     80'h40_E800_80_0000_0C88_2F2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a478_1 ( .OUT(na478_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1349_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a478_2 ( .OUT(na478_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na478_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a478_4 ( .OUT(na478_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1253_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a478_5 ( .OUT(na478_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na478_2_i) );
// C_///AND/D      x114y93     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a479_4 ( .OUT(na479_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1350_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a479_5 ( .OUT(na479_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na479_2_i) );
// C_///AND/D      x121y84     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a480_4 ( .OUT(na480_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1351_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a480_5 ( .OUT(na480_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na480_2_i) );
// C_///AND/D      x117y83     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a481_4 ( .OUT(na481_2_i), .IN1(1'b1), .IN2(na1352_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a481_5 ( .OUT(na481_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na481_2_i) );
// C_AND/D///      x112y78     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a482_1 ( .OUT(na482_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1353_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a482_2 ( .OUT(na482_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na482_1_i) );
// C_///AND/D      x111y71     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a483_4 ( .OUT(na483_2_i), .IN1(na1354_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a483_5 ( .OUT(na483_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na483_2_i) );
// C_///AND/D      x119y84     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a484_4 ( .OUT(na484_2_i), .IN1(na1355_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a484_5 ( .OUT(na484_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na484_2_i) );
// C_AND/D///      x115y86     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a485_1 ( .OUT(na485_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1356_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a485_2 ( .OUT(na485_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na485_1_i) );
// C_AND/D///      x113y84     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1357_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a486_2 ( .OUT(na486_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na486_1_i) );
// C_AND/D///      x103y108     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a487_1 ( .OUT(na487_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1358_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a487_2 ( .OUT(na487_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na487_1_i) );
// C_///AND/D      x116y96     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a488_4 ( .OUT(na488_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1359_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a488_5 ( .OUT(na488_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na488_2_i) );
// C_///AND/D      x106y106     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a489_4 ( .OUT(na489_2_i), .IN1(1'b1), .IN2(na1360_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a489_5 ( .OUT(na489_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na489_2_i) );
// C_AND/D//AND/D      x118y91     80'h40_E800_80_0000_0C88_3C3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a490_1 ( .OUT(na490_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1361_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a490_2 ( .OUT(na490_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na490_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a490_4 ( .OUT(na490_2_i), .IN1(1'b1), .IN2(na1265_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a490_5 ( .OUT(na490_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na490_2_i) );
// C_///AND/D      x113y77     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a491_4 ( .OUT(na491_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1362_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a491_5 ( .OUT(na491_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na491_2_i) );
// C_AND/D//AND/D      x110y102     80'h40_E800_80_0000_0C88_4F3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a492_1 ( .OUT(na492_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1363_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a492_2 ( .OUT(na492_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na492_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a492_4 ( .OUT(na492_2_i), .IN1(1'b1), .IN2(na1267_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a492_5 ( .OUT(na492_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na492_2_i) );
// C_AND/D///      x85y108     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_1 ( .OUT(na493_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1124_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a493_2 ( .OUT(na493_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na493_1_i) );
// C_AND/D///      x87y90     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1126_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a495_2 ( .OUT(na495_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na495_1_i) );
// C_AND/D///      x89y76     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a496_1 ( .OUT(na496_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1127_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a496_2 ( .OUT(na496_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na496_1_i) );
// C_///AND/D      x89y73     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a497_4 ( .OUT(na497_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1128_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a497_5 ( .OUT(na497_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na497_2_i) );
// C_///AND/D      x101y63     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a498_4 ( .OUT(na498_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1129_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a498_5 ( .OUT(na498_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na498_2_i) );
// C_///AND/D      x88y64     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a499_4 ( .OUT(na499_2_i), .IN1(1'b1), .IN2(na1130_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a499_5 ( .OUT(na499_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na499_2_i) );
// C_AND/D///      x93y67     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a500_1 ( .OUT(na500_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1131_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a500_2 ( .OUT(na500_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na500_1_i) );
// C_AND/D///      x110y97     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1132_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a501_2 ( .OUT(na501_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na501_1_i) );
// C_AND/D///      x118y78     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1134_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a503_2 ( .OUT(na503_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na503_1_i) );
// C_///AND/D      x119y77     80'h40_E800_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a504_4 ( .OUT(na504_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3011_2), .IN4(na1135_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a504_5 ( .OUT(na504_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na504_2_i) );
// C_///AND/D      x118y70     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a505_4 ( .OUT(na505_2_i), .IN1(1'b1), .IN2(na1136_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a505_5 ( .OUT(na505_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na505_2_i) );
// C_///AND/D      x115y64     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a506_4 ( .OUT(na506_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1137_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a506_5 ( .OUT(na506_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na506_2_i) );
// C_AND/D///      x111y66     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a507_1 ( .OUT(na507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1138_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a507_2 ( .OUT(na507_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na507_1_i) );
// C_AND/D///      x114y68     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a508_1 ( .OUT(na508_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1139_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a508_2 ( .OUT(na508_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na508_1_i) );
// C_AND/D///      x121y85     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a509_1 ( .OUT(na509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1140_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a509_2 ( .OUT(na509_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na509_1_i) );
// C_///AND/D      x115y80     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a510_4 ( .OUT(na510_2_i), .IN1(1'b1), .IN2(na1141_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a510_5 ( .OUT(na510_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na510_2_i) );
// C_AND/D///      x100y110     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a511_1 ( .OUT(na511_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a511_2 ( .OUT(na511_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na511_1_i) );
// C_///AND/D      x114y101     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a512_4 ( .OUT(na512_2_i), .IN1(1'b1), .IN2(na1143_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a512_5 ( .OUT(na512_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na512_2_i) );
// C_///AND/D      x106y111     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a513_4 ( .OUT(na513_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1144_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a513_5 ( .OUT(na513_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na513_2_i) );
// C_///AND/D      x117y70     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a515_4 ( .OUT(na515_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1146_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a515_5 ( .OUT(na515_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na515_2_i) );
// C_AND/D///      x96y85     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a517_1 ( .OUT(na517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1115_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a517_2 ( .OUT(na517_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na517_1_i) );
// C_AND/D///      x101y107     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a518_1 ( .OUT(na518_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1116_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a518_2 ( .OUT(na518_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na518_1_i) );
// C_AND/D///      x102y106     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a519_1 ( .OUT(na519_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1117_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a519_2 ( .OUT(na519_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na519_1_i) );
// C_///AND/D      x112y96     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a520_4 ( .OUT(na520_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1118_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a520_5 ( .OUT(na520_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na520_2_i) );
// C_///AND/D      x121y85     80'h40_E800_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a521_4 ( .OUT(na521_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3011_2), .IN4(na1120_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a521_5 ( .OUT(na521_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na521_2_i) );
// C_///AND/D      x114y68     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a522_4 ( .OUT(na522_2_i), .IN1(1'b1), .IN2(na1121_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a522_5 ( .OUT(na522_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na522_2_i) );
// C_AND/D///      x110y66     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1122_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a523_2 ( .OUT(na523_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na523_1_i) );
// C_AND/D///      x112y72     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a524_1 ( .OUT(na524_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1123_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a524_2 ( .OUT(na524_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na524_1_i) );
// C_AND/D///      x88y110     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1148_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a525_2 ( .OUT(na525_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na525_1_i) );
// C_///AND/D      x86y109     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a526_4 ( .OUT(na526_2_i), .IN1(1'b1), .IN2(na1149_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a526_5 ( .OUT(na526_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na526_2_i) );
// C_///AND/D      x85y94     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a527_4 ( .OUT(na527_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1150_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a527_5 ( .OUT(na527_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na527_2_i) );
// C_///AND/D      x92y76     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a528_4 ( .OUT(na528_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1151_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a528_5 ( .OUT(na528_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na528_2_i) );
// C_AND/D///      x92y66     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a529_1 ( .OUT(na529_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1152_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a529_2 ( .OUT(na529_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na529_1_i) );
// C_AND/D///      x109y63     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a530_1 ( .OUT(na530_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1153_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a530_2 ( .OUT(na530_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na530_1_i) );
// C_AND/D///      x90y63     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a531_1 ( .OUT(na531_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1154_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a531_2 ( .OUT(na531_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na531_1_i) );
// C_///AND/D      x96y66     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a532_4 ( .OUT(na532_2_i), .IN1(1'b1), .IN2(na1155_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a532_5 ( .OUT(na532_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na532_2_i) );
// C_///AND/D      x109y98     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a533_4 ( .OUT(na533_2_i), .IN1(1'b1), .IN2(na1156_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a533_5 ( .OUT(na533_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na533_2_i) );
// C_///AND/D      x108y106     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a534_4 ( .OUT(na534_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1157_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a534_5 ( .OUT(na534_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na534_2_i) );
// C_AND/D///      x121y81     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a535_1 ( .OUT(na535_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1158_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a535_2 ( .OUT(na535_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na535_1_i) );
// C_///AND/D      x118y77     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a536_4 ( .OUT(na536_2_i), .IN1(1'b1), .IN2(na1159_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a536_5 ( .OUT(na536_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na536_2_i) );
// C_AND/D///      x119y69     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a537_1 ( .OUT(na537_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1160_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a537_2 ( .OUT(na537_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na537_1_i) );
// C_///AND/D      x114y65     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a538_4 ( .OUT(na538_2_i), .IN1(1'b1), .IN2(na1161_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a538_5 ( .OUT(na538_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na538_2_i) );
// C_///AND/D      x115y71     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a539_4 ( .OUT(na539_2_i), .IN1(1'b1), .IN2(na1162_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a539_5 ( .OUT(na539_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na539_2_i) );
// C_AND/D///      x115y70     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a540_1 ( .OUT(na540_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1163_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a540_2 ( .OUT(na540_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na540_1_i) );
// C_AND/D///      x119y81     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a541_1 ( .OUT(na541_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1164_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a541_2 ( .OUT(na541_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na541_1_i) );
// C_///AND/D      x118y75     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a542_4 ( .OUT(na542_2_i), .IN1(1'b1), .IN2(na1165_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a542_5 ( .OUT(na542_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na542_2_i) );
// C_///AND/D      x101y108     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a543_4 ( .OUT(na543_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1166_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a543_5 ( .OUT(na543_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na543_2_i) );
// C_///AND/D      x120y100     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a544_4 ( .OUT(na544_2_i), .IN1(1'b1), .IN2(na1167_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a544_5 ( .OUT(na544_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na544_2_i) );
// C_AND/D///      x107y107     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a545_1 ( .OUT(na545_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1168_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a545_2 ( .OUT(na545_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na545_1_i) );
// C_AND/D///      x120y90     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a546_1 ( .OUT(na546_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1169_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a546_2 ( .OUT(na546_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na546_1_i) );
// C_AND/D///      x118y69     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a547_1 ( .OUT(na547_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1170_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a547_2 ( .OUT(na547_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na547_1_i) );
// C_///AND/D      x111y108     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a548_4 ( .OUT(na548_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1171_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a548_5 ( .OUT(na548_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na548_2_i) );
// C_///AND/D      x96y86     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a549_4 ( .OUT(na549_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1172_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a549_5 ( .OUT(na549_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na549_2_i) );
// C_///AND/D      x103y106     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a550_4 ( .OUT(na550_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1173_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a550_5 ( .OUT(na550_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na550_2_i) );
// C_AND/D///      x100y102     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a551_1 ( .OUT(na551_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1174_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a551_2 ( .OUT(na551_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na551_1_i) );
// C_AND/D///      x115y92     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a552_1 ( .OUT(na552_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1175_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a552_2 ( .OUT(na552_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na552_1_i) );
// C_AND/D///      x118y81     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a553_1 ( .OUT(na553_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1176_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a553_2 ( .OUT(na553_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na553_1_i) );
// C_///AND/D      x117y65     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a554_4 ( .OUT(na554_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1177_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a554_5 ( .OUT(na554_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na554_2_i) );
// C_///AND/D      x105y66     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a555_4 ( .OUT(na555_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1178_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a555_5 ( .OUT(na555_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na555_2_i) );
// C_///AND/D      x111y68     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a556_4 ( .OUT(na556_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1179_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a556_5 ( .OUT(na556_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na556_2_i) );
// C_AND/D///      x89y107     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a557_1 ( .OUT(na557_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1180_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a557_2 ( .OUT(na557_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na557_1_i) );
// C_///AND/D      x85y108     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a558_4 ( .OUT(na558_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1181_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a558_5 ( .OUT(na558_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na558_2_i) );
// C_AND/D///      x86y93     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a559_1 ( .OUT(na559_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1182_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a559_2 ( .OUT(na559_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na559_1_i) );
// C_AND/D///      x90y77     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a560_1 ( .OUT(na560_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1183_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a560_2 ( .OUT(na560_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na560_1_i) );
// C_AND/D///      x89y68     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a561_1 ( .OUT(na561_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1184_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a561_2 ( .OUT(na561_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na561_1_i) );
// C_///AND/D      x106y64     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a562_4 ( .OUT(na562_2_i), .IN1(1'b1), .IN2(na1185_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a562_5 ( .OUT(na562_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na562_2_i) );
// C_///AND/D      x86y64     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a563_4 ( .OUT(na563_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1186_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a563_5 ( .OUT(na563_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na563_2_i) );
// C_///AND/D      x94y68     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a564_4 ( .OUT(na564_2_i), .IN1(1'b1), .IN2(na1187_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a564_5 ( .OUT(na564_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na564_2_i) );
// C_AND/D///      x110y100     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a565_1 ( .OUT(na565_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1188_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a565_2 ( .OUT(na565_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na565_1_i) );
// C_AND/D///      x107y112     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a566_1 ( .OUT(na566_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1189_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a566_2 ( .OUT(na566_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na566_1_i) );
// C_AND/D///      x118y84     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1190_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a567_2 ( .OUT(na567_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na567_1_i) );
// C_AND/D///      x121y78     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a568_1 ( .OUT(na568_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1191_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a568_2 ( .OUT(na568_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na568_1_i) );
// C_AND/D///      x116y73     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_1 ( .OUT(na569_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1192_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a569_2 ( .OUT(na569_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na569_1_i) );
// C_AND/D///      x113y65     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a570_1 ( .OUT(na570_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1193_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a570_2 ( .OUT(na570_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na570_1_i) );
// C_AND/D///      x112y70     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a571_1 ( .OUT(na571_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1194_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a571_2 ( .OUT(na571_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na571_1_i) );
// C_///AND/D      x113y70     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a572_4 ( .OUT(na572_2_i), .IN1(1'b1), .IN2(na1195_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a572_5 ( .OUT(na572_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na572_2_i) );
// C_AND/D///      x117y84     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a573_1 ( .OUT(na573_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1196_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a573_2 ( .OUT(na573_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na573_1_i) );
// C_///AND/D      x114y78     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a574_4 ( .OUT(na574_2_i), .IN1(na1197_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a574_5 ( .OUT(na574_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na574_2_i) );
// C_AND/D///      x102y109     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a575_1 ( .OUT(na575_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1198_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a575_2 ( .OUT(na575_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na575_1_i) );
// C_///AND/D      x114y97     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a576_4 ( .OUT(na576_2_i), .IN1(1'b1), .IN2(na1199_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a576_5 ( .OUT(na576_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na576_2_i) );
// C_AND/D///      x103y106     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_1 ( .OUT(na577_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1200_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a577_2 ( .OUT(na577_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na577_1_i) );
// C_///AND/D      x121y94     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a578_4 ( .OUT(na578_2_i), .IN1(1'b1), .IN2(~na3013_2), .IN3(1'b1), .IN4(na1201_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a578_5 ( .OUT(na578_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na578_2_i) );
// C_AND/D///      x115y72     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_1 ( .OUT(na579_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1202_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a579_2 ( .OUT(na579_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na579_1_i) );
// C_///AND/D      x108y108     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a580_4 ( .OUT(na580_2_i), .IN1(1'b1), .IN2(na1203_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a580_5 ( .OUT(na580_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na580_2_i) );
// C_AND/D///      x95y88     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_1 ( .OUT(na581_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1204_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a581_2 ( .OUT(na581_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na581_1_i) );
// C_///AND/D      x95y110     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a582_4 ( .OUT(na582_2_i), .IN1(1'b1), .IN2(na1205_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a582_5 ( .OUT(na582_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na582_2_i) );
// C_AND/D///      x97y106     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_1 ( .OUT(na583_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1206_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a583_2 ( .OUT(na583_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na583_1_i) );
// C_///AND/D      x114y98     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a584_4 ( .OUT(na584_2_i), .IN1(na1207_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a584_5 ( .OUT(na584_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na584_2_i) );
// C_AND/D///      x115y82     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_1 ( .OUT(na585_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1208_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a585_2 ( .OUT(na585_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na585_1_i) );
// C_///AND/D      x118y65     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a586_4 ( .OUT(na586_2_i), .IN1(1'b1), .IN2(~na3013_2), .IN3(1'b1), .IN4(na1209_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a586_5 ( .OUT(na586_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na586_2_i) );
// C_AND/D///      x105y66     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_1 ( .OUT(na587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1210_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a587_2 ( .OUT(na587_1), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na587_1_i) );
// C_///AND/D      x106y68     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a588_4 ( .OUT(na588_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1211_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a588_5 ( .OUT(na588_2), .CLK(1'b0), .EN(na1111_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na588_2_i) );
// C_AND/D///      x87y107     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a589_1 ( .OUT(na589_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1244_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a589_2 ( .OUT(na589_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na589_1_i) );
// C_///AND/D      x86y90     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a591_4 ( .OUT(na591_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1246_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a591_5 ( .OUT(na591_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na591_2_i) );
// C_AND/D///      x87y77     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a592_1 ( .OUT(na592_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1247_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a592_2 ( .OUT(na592_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na592_1_i) );
// C_///AND/D      x91y68     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a593_4 ( .OUT(na593_2_i), .IN1(1'b1), .IN2(na1248_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a593_5 ( .OUT(na593_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na593_2_i) );
// C_AND/D///      x99y64     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_1 ( .OUT(na594_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1249_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a594_2 ( .OUT(na594_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na594_1_i) );
// C_///AND/D      x92y63     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a595_4 ( .OUT(na595_2_i), .IN1(1'b1), .IN2(na1250_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a595_5 ( .OUT(na595_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na595_2_i) );
// C_AND/D///      x92y67     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a596_1 ( .OUT(na596_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1251_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a596_2 ( .OUT(na596_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na596_1_i) );
// C_///AND/D      x119y93     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a597_4 ( .OUT(na597_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1252_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a597_5 ( .OUT(na597_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na597_2_i) );
// C_AND/D///      x120y81     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a599_1 ( .OUT(na599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1254_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a599_2 ( .OUT(na599_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na599_1_i) );
// C_///AND/D      x118y71     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a600_4 ( .OUT(na600_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1255_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a600_5 ( .OUT(na600_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na600_2_i) );
// C_AND/D///      x118y71     80'h40_E800_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a601_1 ( .OUT(na601_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1256_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a601_2 ( .OUT(na601_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na601_1_i) );
// C_///AND/D      x115y65     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a602_4 ( .OUT(na602_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1257_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a602_5 ( .OUT(na602_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na602_2_i) );
// C_AND/D///      x112y66     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a603_1 ( .OUT(na603_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1258_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a603_2 ( .OUT(na603_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na603_1_i) );
// C_///AND/D      x116y65     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a604_4 ( .OUT(na604_2_i), .IN1(na1259_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a604_5 ( .OUT(na604_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na604_2_i) );
// C_AND/D///      x119y84     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a605_1 ( .OUT(na605_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1260_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a605_2 ( .OUT(na605_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na605_1_i) );
// C_///AND/D      x114y76     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a606_4 ( .OUT(na606_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1261_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a606_5 ( .OUT(na606_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na606_2_i) );
// C_AND/D///      x101y110     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a607_1 ( .OUT(na607_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1262_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a607_2 ( .OUT(na607_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na607_1_i) );
// C_///AND/D      x115y97     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a608_4 ( .OUT(na608_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1263_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a608_5 ( .OUT(na608_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na608_2_i) );
// C_AND/D///      x107y110     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a609_1 ( .OUT(na609_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1264_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a609_2 ( .OUT(na609_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na609_1_i) );
// C_///AND/D      x116y72     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a611_4 ( .OUT(na611_2_i), .IN1(1'b1), .IN2(na1266_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a611_5 ( .OUT(na611_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na611_2_i) );
// C_AND/D///      x88y103     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a615_1 ( .OUT(na615_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1270_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a615_2 ( .OUT(na615_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na615_1_i) );
// C_///AND/D      x109y102     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a616_4 ( .OUT(na616_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1271_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a616_5 ( .OUT(na616_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na616_2_i) );
// C_AND/D///      x113y90     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a617_1 ( .OUT(na617_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1272_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a617_2 ( .OUT(na617_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na617_1_i) );
// C_///AND/D      x112y67     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a618_4 ( .OUT(na618_2_i), .IN1(na1273_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a618_5 ( .OUT(na618_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na618_2_i) );
// C_AND/D///      x92y109     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a621_1 ( .OUT(na621_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1276_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a621_2 ( .OUT(na621_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na621_1_i) );
// C_///AND/D      x88y109     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a622_4 ( .OUT(na622_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1277_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a622_5 ( .OUT(na622_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na622_2_i) );
// C_AND/D///      x87y93     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a623_1 ( .OUT(na623_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1278_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a623_2 ( .OUT(na623_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na623_1_i) );
// C_///AND/D      x89y77     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a624_4 ( .OUT(na624_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1279_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a624_5 ( .OUT(na624_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na624_2_i) );
// C_///AND/D      x94y66     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a625_4 ( .OUT(na625_2_i), .IN1(na1280_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a625_5 ( .OUT(na625_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na625_2_i) );
// C_///AND/D      x107y63     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a626_4 ( .OUT(na626_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1281_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a626_5 ( .OUT(na626_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na626_2_i) );
// C_AND/D///      x94y64     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a627_1 ( .OUT(na627_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1282_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a627_2 ( .OUT(na627_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na627_1_i) );
// C_AND/D///      x95y68     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a628_1 ( .OUT(na628_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1283_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a628_2 ( .OUT(na628_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na628_1_i) );
// C_///AND/D      x119y95     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a629_4 ( .OUT(na629_2_i), .IN1(1'b1), .IN2(na1284_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a629_5 ( .OUT(na629_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na629_2_i) );
// C_AND/D///      x108y105     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a630_1 ( .OUT(na630_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1285_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a630_2 ( .OUT(na630_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na630_1_i) );
// C_AND/D///      x123y85     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a631_1 ( .OUT(na631_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1286_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a631_2 ( .OUT(na631_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na631_1_i) );
// C_AND/D///      x118y74     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a632_1 ( .OUT(na632_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1287_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a632_2 ( .OUT(na632_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na632_1_i) );
// C_///AND/D      x122y71     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a633_4 ( .OUT(na633_2_i), .IN1(na1288_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a633_5 ( .OUT(na633_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na633_2_i) );
// C_AND/D///      x116y68     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a634_1 ( .OUT(na634_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1289_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a634_2 ( .OUT(na634_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na634_1_i) );
// C_///AND/D      x113y72     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a635_4 ( .OUT(na635_2_i), .IN1(1'b1), .IN2(~na3013_2), .IN3(1'b1), .IN4(na1290_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a635_5 ( .OUT(na635_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na635_2_i) );
// C_AND/D///      x116y72     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a636_1 ( .OUT(na636_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1291_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a636_2 ( .OUT(na636_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na636_1_i) );
// C_///AND/D      x120y82     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a637_4 ( .OUT(na637_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1292_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a637_5 ( .OUT(na637_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na637_2_i) );
// C_AND/D///      x114y76     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a638_1 ( .OUT(na638_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1293_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a638_2 ( .OUT(na638_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na638_1_i) );
// C_///AND/D      x103y107     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a639_4 ( .OUT(na639_2_i), .IN1(1'b1), .IN2(~na3013_2), .IN3(1'b1), .IN4(na1294_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a639_5 ( .OUT(na639_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na639_2_i) );
// C_AND/D///      x115y97     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a640_1 ( .OUT(na640_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1295_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a640_2 ( .OUT(na640_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na640_1_i) );
// C_///AND/D      x104y107     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a641_4 ( .OUT(na641_2_i), .IN1(1'b1), .IN2(na1296_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a641_5 ( .OUT(na641_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na641_2_i) );
// C_AND/D///      x118y90     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a642_1 ( .OUT(na642_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1297_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a642_2 ( .OUT(na642_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na642_1_i) );
// C_///AND/D      x116y68     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a643_4 ( .OUT(na643_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1298_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a643_5 ( .OUT(na643_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na643_2_i) );
// C_AND/D///      x110y103     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a644_1 ( .OUT(na644_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1299_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a644_2 ( .OUT(na644_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na644_1_i) );
// C_///AND/D      x86y101     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a645_4 ( .OUT(na645_2_i), .IN1(na1300_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a645_5 ( .OUT(na645_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na645_2_i) );
// C_AND/D///      x95y109     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a646_1 ( .OUT(na646_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1301_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a646_2 ( .OUT(na646_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na646_1_i) );
// C_///AND/D      x94y107     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a647_4 ( .OUT(na647_2_i), .IN1(1'b1), .IN2(na1302_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a647_5 ( .OUT(na647_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na647_2_i) );
// C_AND/D///      x105y97     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a648_1 ( .OUT(na648_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1303_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a648_2 ( .OUT(na648_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na648_1_i) );
// C_///AND/D      x112y90     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a649_4 ( .OUT(na649_2_i), .IN1(na1304_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a649_5 ( .OUT(na649_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na649_2_i) );
// C_AND/D///      x115y66     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a650_1 ( .OUT(na650_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1305_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a650_2 ( .OUT(na650_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na650_1_i) );
// C_///AND/D      x103y65     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a651_4 ( .OUT(na651_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1306_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a651_5 ( .OUT(na651_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na651_2_i) );
// C_AND/D///      x108y70     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a652_1 ( .OUT(na652_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1307_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a652_2 ( .OUT(na652_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na652_1_i) );
// C_///AND/D      x88y108     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a653_4 ( .OUT(na653_2_i), .IN1(1'b1), .IN2(na1308_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a653_5 ( .OUT(na653_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na653_2_i) );
// C_AND/D///      x85y107     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a654_1 ( .OUT(na654_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1309_1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a654_2 ( .OUT(na654_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na654_1_i) );
// C_///AND/D      x87y96     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a655_4 ( .OUT(na655_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1310_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a655_5 ( .OUT(na655_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na655_2_i) );
// C_AND/D///      x90y79     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a656_1 ( .OUT(na656_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1311_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a656_2 ( .OUT(na656_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na656_1_i) );
// C_///AND/D      x88y63     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a657_4 ( .OUT(na657_2_i), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(na1312_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a657_5 ( .OUT(na657_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na657_2_i) );
// C_AND/D///      x108y64     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a658_1 ( .OUT(na658_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1313_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a658_2 ( .OUT(na658_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na658_1_i) );
// C_///AND/D      x96y63     80'h40_E800_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a659_4 ( .OUT(na659_2_i), .IN1(1'b1), .IN2(~na3013_2), .IN3(1'b1), .IN4(na1314_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a659_5 ( .OUT(na659_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na659_2_i) );
// C_AND/D///      x95y66     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a660_1 ( .OUT(na660_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1315_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a660_2 ( .OUT(na660_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na660_1_i) );
// C_///AND/D      x118y96     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a661_4 ( .OUT(na661_2_i), .IN1(1'b1), .IN2(na1316_1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a661_5 ( .OUT(na661_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na661_2_i) );
// C_AND/D///      x107y106     80'h40_E800_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a662_1 ( .OUT(na662_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3011_2), .IN8(na1317_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a662_2 ( .OUT(na662_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na662_1_i) );
// C_///AND/D      x118y90     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a663_4 ( .OUT(na663_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1318_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a663_5 ( .OUT(na663_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na663_2_i) );
// C_AND/D///      x117y76     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a664_1 ( .OUT(na664_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1319_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a664_2 ( .OUT(na664_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na664_1_i) );
// C_///AND/D      x117y76     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a665_4 ( .OUT(na665_2_i), .IN1(1'b1), .IN2(na1320_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a665_5 ( .OUT(na665_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na665_2_i) );
// C_AND/D///      x115y69     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a666_1 ( .OUT(na666_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1321_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a666_2 ( .OUT(na666_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na666_1_i) );
// C_///AND/D      x114y71     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a667_4 ( .OUT(na667_2_i), .IN1(1'b1), .IN2(na1322_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a667_5 ( .OUT(na667_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na667_2_i) );
// C_AND/D///      x115y73     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a668_1 ( .OUT(na668_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1323_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a668_2 ( .OUT(na668_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na668_1_i) );
// C_///AND/D      x121y83     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a669_4 ( .OUT(na669_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1324_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a669_5 ( .OUT(na669_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na669_2_i) );
// C_AND/D///      x113y78     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a670_1 ( .OUT(na670_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1325_2), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a670_2 ( .OUT(na670_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na670_1_i) );
// C_///AND/D      x104y111     80'h40_E800_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a671_4 ( .OUT(na671_2_i), .IN1(1'b1), .IN2(na1326_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a671_5 ( .OUT(na671_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na671_2_i) );
// C_AND/D///      x113y100     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a672_1 ( .OUT(na672_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1327_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a672_2 ( .OUT(na672_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na672_1_i) );
// C_///AND/D      x105y109     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a673_4 ( .OUT(na673_2_i), .IN1(na1328_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a673_5 ( .OUT(na673_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na673_2_i) );
// C_AND/D///      x117y90     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a674_1 ( .OUT(na674_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1329_1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a674_2 ( .OUT(na674_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na674_1_i) );
// C_///AND/D      x116y71     80'h40_E800_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a675_4 ( .OUT(na675_2_i), .IN1(na1330_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a675_5 ( .OUT(na675_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na675_2_i) );
// C_AND/D///      x109y102     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a676_1 ( .OUT(na676_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1331_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a676_2 ( .OUT(na676_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na676_1_i) );
// C_///AND/D      x87y102     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a677_4 ( .OUT(na677_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1332_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a677_5 ( .OUT(na677_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na677_2_i) );
// C_AND/D///      x94y109     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a678_1 ( .OUT(na678_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1333_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a678_2 ( .OUT(na678_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na678_1_i) );
// C_///AND/D      x91y106     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a679_4 ( .OUT(na679_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1334_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a679_5 ( .OUT(na679_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na679_2_i) );
// C_AND/D///      x105y98     80'h40_E800_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a680_1 ( .OUT(na680_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3013_2), .IN7(1'b1), .IN8(na1335_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a680_2 ( .OUT(na680_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na680_1_i) );
// C_///AND/D      x108y83     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a681_4 ( .OUT(na681_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1336_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a681_5 ( .OUT(na681_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na681_2_i) );
// C_AND/D///      x112y67     80'h40_E800_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a682_1 ( .OUT(na682_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1337_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a682_2 ( .OUT(na682_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na682_1_i) );
// C_///AND/D      x104y65     80'h40_E800_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a683_4 ( .OUT(na683_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1338_2), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a683_5 ( .OUT(na683_2), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na683_2_i) );
// C_AND/D///      x108y67     80'h40_E800_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a684_1 ( .OUT(na684_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1339_2), .IN7(1'b1), .IN8(~na429_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a684_2 ( .OUT(na684_1), .CLK(1'b0), .EN(na1112_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na684_1_i) );
// C_AND/D//AND/D      x116y93     80'h40_E800_80_0000_0C88_F4A3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3061_2), .IN6(na686_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a685_2 ( .OUT(na685_1), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na685_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a685_4 ( .OUT(na685_2_i), .IN1(1'b1), .IN2(~na686_1), .IN3(na685_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a685_5 ( .OUT(na685_2), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na685_2_i) );
// C_AND////D      x113y80     80'h40_E818_00_0000_0888_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a686_1 ( .OUT(na686_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1087_2), .IN6(na2923_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a686_5 ( .OUT(na686_2), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na686_1) );
// C_AND/D//AND/D      x117y79     80'h40_E800_80_0000_0C88_A3F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a688_1 ( .OUT(na688_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na686_1), .IN7(na685_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a688_2 ( .OUT(na688_1), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na688_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a688_4 ( .OUT(na688_2_i), .IN1(na688_1), .IN2(~na686_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a688_5 ( .OUT(na688_2), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na688_2_i) );
// C_AND/D//AND/D      x118y67     80'h40_E800_80_0000_0C88_F2A3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a690_1 ( .OUT(na690_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na688_2), .IN6(~na686_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a690_2 ( .OUT(na690_1), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na690_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a690_4 ( .OUT(na690_2_i), .IN1(1'b1), .IN2(~na686_1), .IN3(na690_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a690_5 ( .OUT(na690_2), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na690_2_i) );
// C_///AND/D      x116y70     80'h40_E800_80_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a692_4 ( .OUT(na692_2_i), .IN1(1'b1), .IN2(~na686_1), .IN3(na690_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a692_5 ( .OUT(na692_2), .CLK(1'b0), .EN(na1099_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na692_2_i) );
// C_XOR////D      x122y79     80'h40_E818_00_0000_0666_9AA9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a693_1 ( .OUT(na693_1), .IN1(~na721_1), .IN2(na718_1), .IN3(na732_1), .IN4(1'b0), .IN5(na695_2), .IN6(1'b0), .IN7(~na723_1),
                     .IN8(na3081_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a693_5 ( .OUT(na693_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na693_1) );
// C_///ANDXOR/      x121y77     80'h00_0060_00_0000_0C06_FFD7
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a695_4 ( .OUT(na695_2), .IN1(na696_1), .IN2(na3067_2), .IN3(na717_1), .IN4(~na702_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y71     80'h00_0018_00_0040_0AF8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a696_1 ( .OUT(na696_1), .IN1(na1458_1), .IN2(1'b1), .IN3(~na709_1), .IN4(1'b1), .IN5(na3062_2), .IN6(na713_1), .IN7(na2668_2),
                     .IN8(~na697_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y74     80'h00_0018_00_0040_0AF9_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a697_1 ( .OUT(na697_1), .IN1(na703_2), .IN2(1'b1), .IN3(1'b1), .IN4(na700_2), .IN5(~na703_1), .IN6(na3065_2), .IN7(na3071_2),
                     .IN8(~na700_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y84     80'h00_0018_00_0040_0A73_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a699_1 ( .OUT(na699_1), .IN1(1'b1), .IN2(na704_2), .IN3(1'b1), .IN4(na700_1), .IN5(~na1045_1), .IN6(~na704_1), .IN7(na2670_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x126y80     80'h00_0078_00_0000_0C66_3A60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a700_1 ( .OUT(na700_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1043_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1039_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a700_4 ( .OUT(na700_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2669_1), .IN4(na699_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x124y80     80'h00_0078_00_0000_0C66_6696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1045_1), .IN6(~na1049_1), .IN7(na1041_1),
                     .IN8(na1039_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a702_4 ( .OUT(na702_2), .IN1(na1043_1), .IN2(na1049_1), .IN3(na1037_1), .IN4(~na1047_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x123y77     80'h00_0078_00_0000_0C66_AC09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na704_1), .IN7(na1035_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a703_4 ( .OUT(na703_2), .IN1(~na1045_1), .IN2(na1049_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x123y82     80'h00_0078_00_0000_0C66_9A5C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a704_1 ( .OUT(na704_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1043_1), .IN6(1'b0), .IN7(na3138_2), .IN8(~na1047_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a704_4 ( .OUT(na704_2), .IN1(1'b0), .IN2(na1049_1), .IN3(~na1037_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x124y83     80'h00_0078_00_0000_0C66_C560
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a706_1 ( .OUT(na706_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na703_1), .IN6(1'b0), .IN7(1'b0), .IN8(na700_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a706_4 ( .OUT(na706_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1037_1), .IN4(na1039_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y88     80'h00_0018_00_0040_0A64_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1), .IN1(~na3137_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3139_2), .IN5(1'b0), .IN6(na1049_1), .IN7(~na3140_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y77     80'h00_0018_00_0000_0666_A665
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1), .IN1(~na1045_1), .IN2(1'b0), .IN3(na2671_2), .IN4(na702_1), .IN5(~na711_1), .IN6(~na3135_2), .IN7(na2671_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y83     80'h00_0018_00_0040_0AD9_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1), .IN1(1'b1), .IN2(na704_1), .IN3(1'b1), .IN4(~na700_1), .IN5(~na3134_2), .IN6(1'b0), .IN7(na2672_1),
                     .IN8(~na702_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x123y78     80'h00_0018_00_0000_0666_D5BE
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a713_1 ( .OUT(na713_1), .IN1(~na3073_2), .IN2(~na704_1), .IN3(~na706_1), .IN4(na702_1), .IN5(na716_1), .IN6(1'b1), .IN7(na706_2),
                     .IN8(~na702_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x123y81     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a716_1 ( .OUT(na716_1), .IN1(~na703_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1043_1), .IN6(na2677_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y71     80'h00_0018_00_0040_0AF8_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a717_1 ( .OUT(na717_1), .IN1(1'b1), .IN2(na713_1), .IN3(na709_1), .IN4(1'b1), .IN5(na1458_1), .IN6(na2678_2), .IN7(na3063_2),
                     .IN8(~na697_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y76     80'h00_0018_00_0040_0ABC_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a718_1 ( .OUT(na718_1), .IN1(1'b1), .IN2(~na720_1), .IN3(na719_1), .IN4(1'b1), .IN5(na703_2), .IN6(na704_1), .IN7(1'b1),
                     .IN8(~na3086_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y69     80'h00_0018_00_0040_0AF3_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1), .IN1(1'b1), .IN2(na713_1), .IN3(1'b1), .IN4(~na3163_2), .IN5(~na2680_1), .IN6(~na3075_2), .IN7(na3184_2),
                     .IN8(na697_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y70     80'h00_0018_00_0040_0AF5_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a720_1 ( .OUT(na720_1), .IN1(na1458_1), .IN2(1'b1), .IN3(1'b1), .IN4(na697_1), .IN5(~na3076_2), .IN6(na713_1), .IN7(~na709_1),
                     .IN8(na2682_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y83     80'h00_0018_00_0040_0AED_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1), .IN1(na696_1), .IN2(1'b1), .IN3(~na719_1), .IN4(1'b1), .IN5(1'b1), .IN6(na722_1), .IN7(~na1035_1),
                     .IN8(~na729_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y68     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a722_1 ( .OUT(na722_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na703_2), .IN6(1'b0), .IN7(1'b0), .IN8(na700_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y77     80'h00_0018_00_0040_0AE7_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1), .IN1(1'b1), .IN2(~na720_1), .IN3(na717_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3080_2), .IN7(~na724_1),
                     .IN8(na2684_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y63     80'h00_0018_00_0000_0C66_3C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a724_1 ( .OUT(na724_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na704_2), .IN7(1'b0), .IN8(~na702_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y73     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a725_4 ( .OUT(na725_2), .IN1(1'b0), .IN2(na3068_2), .IN3(~na1037_1), .IN4(na1039_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y77     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a726_1 ( .OUT(na726_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na727_1), .IN8(na730_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y67     80'h00_0018_00_0040_0A72_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1), .IN1(na3077_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3078_2), .IN5(na2685_1), .IN6(~na3186_2), .IN7(na724_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x122y76     80'h00_0078_00_0000_0C66_60A3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a729_1 ( .OUT(na729_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1041_1), .IN8(na1039_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a729_4 ( .OUT(na729_2), .IN1(1'b0), .IN2(~na722_1), .IN3(na1035_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y72     80'h00_0018_00_0040_0ADB_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a730_1 ( .OUT(na730_1), .IN1(~na696_1), .IN2(1'b1), .IN3(na717_1), .IN4(1'b1), .IN5(~na725_2), .IN6(1'b1), .IN7(na2686_2),
                     .IN8(~na729_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y71     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a732_1 ( .OUT(na732_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na734_1), .IN6(na733_1), .IN7(~na3085_2), .IN8(na736_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y72     80'h00_0018_00_0040_0A79_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a733_1 ( .OUT(na733_1), .IN1(~na696_1), .IN2(1'b1), .IN3(na719_1), .IN4(1'b1), .IN5(~na737_1), .IN6(na704_1), .IN7(na3072_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y73     80'h00_0018_00_0040_0AB5_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a734_1 ( .OUT(na734_1), .IN1(1'b1), .IN2(~na720_1), .IN3(~na717_1), .IN4(1'b1), .IN5(~na3066_2), .IN6(na2688_1), .IN7(1'b1),
                     .IN8(na702_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y82     80'h00_0018_00_0040_0AE9_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a735_1 ( .OUT(na735_1), .IN1(1'b1), .IN2(~na720_1), .IN3(~na719_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2688_1), .IN7(na3070_2),
                     .IN8(~na702_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y80     80'h00_0018_00_0040_0ADB_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a736_1 ( .OUT(na736_1), .IN1(~na696_1), .IN2(1'b1), .IN3(na717_1), .IN4(1'b1), .IN5(~na737_1), .IN6(1'b1), .IN7(na2690_2),
                     .IN8(~na729_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y75     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na703_2), .IN6(na704_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x115y84     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a738_1 ( .OUT(na738_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na2691_1), .IN6(1'b0), .IN7(na693_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a738_2 ( .OUT(na738_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na738_1_i) );
// C_XOR////D      x117y91     80'h40_E818_00_0000_0666_696A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1), .IN1(na726_1), .IN2(1'b0), .IN3(~na744_1), .IN4(~na741_2), .IN5(na721_1), .IN6(~na735_1), .IN7(na723_1),
                     .IN8(na736_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a739_5 ( .OUT(na739_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na739_1) );
// C_///XOR/      x124y66     80'h00_0060_00_0000_0C06_FF96
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a741_4 ( .OUT(na741_2), .IN1(na695_2), .IN2(na718_1), .IN3(na3089_2), .IN4(~na742_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y64     80'h00_0018_00_0040_0AB8_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a742_1 ( .OUT(na742_1), .IN1(1'b1), .IN2(~na720_1), .IN3(na719_1), .IN4(1'b1), .IN5(na725_2), .IN6(na3079_2), .IN7(1'b0),
                     .IN8(~na2684_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y64     80'h00_0018_00_0040_0AE7_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a743_1 ( .OUT(na743_1), .IN1(na696_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2693_2), .IN5(1'b1), .IN6(~na3084_2), .IN7(~na717_1),
                     .IN8(na2693_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y65     80'h00_0018_00_0000_0666_56AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a744_1 ( .OUT(na744_1), .IN1(1'b0), .IN2(na733_1), .IN3(na2694_2), .IN4(1'b0), .IN5(na734_1), .IN6(na746_1), .IN7(~na2694_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y64     80'h00_0018_00_0040_0A7C_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a746_1 ( .OUT(na746_1), .IN1(~na696_1), .IN2(1'b1), .IN3(na719_1), .IN4(1'b1), .IN5(na2696_2), .IN6(na722_1), .IN7(~na724_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x105y93     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a747_1 ( .OUT(na747_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na739_1), .IN6(1'b0), .IN7(na2697_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a747_2 ( .OUT(na747_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na747_1_i) );
// C_XOR////D      x115y81     80'h40_E818_00_0000_0666_0ACA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a748_1 ( .OUT(na748_1), .IN1(na749_1), .IN2(1'b0), .IN3(1'b0), .IN4(na752_2), .IN5(na750_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a748_5 ( .OUT(na748_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na748_1) );
// C_XOR////      x121y83     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a749_1 ( .OUT(na749_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na726_1), .IN6(1'b0), .IN7(~na744_1), .IN8(na741_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y79     80'h00_0018_00_0000_0666_9969
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a750_1 ( .OUT(na750_1), .IN1(na695_2), .IN2(~na735_1), .IN3(~na732_1), .IN4(~na741_2), .IN5(~na721_1), .IN6(na718_1), .IN7(~na723_1),
                     .IN8(na736_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x120y84     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a752_4 ( .OUT(na752_2), .IN1(~na695_2), .IN2(~na718_1), .IN3(na732_1), .IN4(na3082_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x105y86     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_1 ( .OUT(na753_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na748_1), .IN6(1'b0), .IN7(na2698_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a753_2 ( .OUT(na753_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na753_1_i) );
// C_XOR////D      x111y75     80'h40_E818_00_0000_0666_C009
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a754_1 ( .OUT(na754_1), .IN1(na750_1), .IN2(~na755_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na752_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a754_5 ( .OUT(na754_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na754_1) );
// C_XOR////      x121y68     80'h00_0018_00_0000_0666_90A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a755_1 ( .OUT(na755_1), .IN1(na758_1), .IN2(na743_1), .IN3(na732_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na757_1),
                     .IN8(na742_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y65     80'h00_0018_00_0040_0A7C_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a757_1 ( .OUT(na757_1), .IN1(1'b1), .IN2(na720_1), .IN3(na719_1), .IN4(1'b1), .IN5(na703_2), .IN6(na2699_1), .IN7(~na3083_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y67     80'h00_0018_00_0040_0AB8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a758_1 ( .OUT(na758_1), .IN1(na696_1), .IN2(1'b1), .IN3(~na717_1), .IN4(1'b1), .IN5(na737_1), .IN6(na2700_2), .IN7(1'b0),
                     .IN8(~na702_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x103y80     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_1 ( .OUT(na759_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na754_1), .IN6(1'b0), .IN7(na2701_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a759_2 ( .OUT(na759_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na759_1_i) );
// C_XOR////D      x108y69     80'h40_E818_00_0000_0666_0C3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a760_1 ( .OUT(na760_1), .IN1(na750_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na761_1), .IN5(1'b0), .IN6(na755_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a760_5 ( .OUT(na760_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na760_1) );
// C_XOR////      x122y66     80'h00_0018_00_0000_0666_66A0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a761_1 ( .OUT(na761_1), .IN1(1'b0), .IN2(1'b0), .IN3(na732_1), .IN4(1'b0), .IN5(na3187_2), .IN6(na746_1), .IN7(na2694_2),
                     .IN8(na741_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x102y77     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a763_1 ( .OUT(na763_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na2702_2), .IN6(1'b0), .IN7(na760_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a763_2 ( .OUT(na763_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na763_1_i) );
// C_XOR////D      x112y61     80'h40_E818_00_0000_0666_0C0A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a764_1 ( .OUT(na764_1), .IN1(na765_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na766_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a764_5 ( .OUT(na764_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na764_1) );
// C_XOR////      x117y63     80'h00_0018_00_0000_0666_9696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1), .IN1(na3088_2), .IN2(na743_1), .IN3(na2694_1), .IN4(~na742_1), .IN5(na758_1), .IN6(na746_1), .IN7(~na757_1),
                     .IN8(na3188_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y64     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a766_1 ( .OUT(na766_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na726_1), .IN6(na743_1), .IN7(na732_1), .IN8(na742_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x104y70     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a768_1 ( .OUT(na768_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na2703_1), .IN6(1'b0), .IN7(na764_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a768_2 ( .OUT(na768_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na768_1_i) );
// C_XOR////D      x107y65     80'h40_E818_00_0000_0666_A005
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a769_1 ( .OUT(na769_1), .IN1(~na765_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na744_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a769_5 ( .OUT(na769_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na769_1) );
// C_MX2b/D///      x100y71     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a770_1 ( .OUT(na770_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na769_1), .IN6(1'b0), .IN7(na2704_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a770_2 ( .OUT(na770_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na770_1_i) );
// C_XOR////D      x107y66     80'h40_E818_00_0000_0666_0C0A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a771_1 ( .OUT(na771_1), .IN1(na765_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na772_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a771_5 ( .OUT(na771_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na771_1) );
// C_///XOR/      x119y64     80'h00_0060_00_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a772_4 ( .OUT(na772_2), .IN1(na726_1), .IN2(na743_1), .IN3(~na744_1), .IN4(~na742_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x102y71     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a773_1 ( .OUT(na773_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b0), .IN6(na771_1), .IN7(1'b0), .IN8(na3195_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a773_2 ( .OUT(na773_1), .CLK(1'b0), .EN(na1096_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na773_1_i) );
// C_XOR////D      x109y100     80'h40_E818_00_0000_0666_A0C0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a774_1 ( .OUT(na774_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na775_1), .IN5(1'b0), .IN6(1'b0), .IN7(na816_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a774_5 ( .OUT(na774_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na774_1) );
// C_XOR////      x120y98     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na814_1), .IN6(na815_1), .IN7(na3092_2), .IN8(na807_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x124y106     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a776_4 ( .OUT(na776_2), .IN1(1'b0), .IN2(na801_1), .IN3(1'b0), .IN4(na777_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y108     80'h00_0018_00_0040_0AE0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1), .IN1(~na778_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2706_2), .IN5(1'b0), .IN6(na2724_2), .IN7(na797_1),
                     .IN8(na2706_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y101     80'h00_0018_00_0040_0AFC_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a778_1 ( .OUT(na778_1), .IN1(na786_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1461_1), .IN5(na2707_2), .IN6(na3197_2), .IN7(~na3196_2),
                     .IN8(~na3100_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y108     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1053_1), .IN8(na1065_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y99     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a780_4 ( .OUT(na780_2), .IN1(na1059_1), .IN2(~na3143_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x124y96     80'h00_0078_00_0000_0C66_6669
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1055_1), .IN6(na1057_1), .IN7(~na1061_1),
                     .IN8(~na1065_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a781_4 ( .OUT(na781_2), .IN1(na1059_1), .IN2(~na1063_1), .IN3(na1053_1), .IN4(na1065_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x122y97     80'h00_0078_00_0000_0C66_9CAA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2716_2), .IN7(na780_2), .IN8(~na1051_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a783_4 ( .OUT(na783_2), .IN1(na1055_1), .IN2(1'b0), .IN3(na1053_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y98     80'h00_0018_00_0040_0A98_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a784_1 ( .OUT(na784_1), .IN1(na1055_1), .IN2(1'b1), .IN3(na1061_1), .IN4(1'b1), .IN5(na3144_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na1065_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x123y97     80'h00_0018_00_0000_0666_D3BE
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a786_1 ( .OUT(na786_1), .IN1(~na3093_2), .IN2(~na2716_2), .IN3(~na783_1), .IN4(na781_1), .IN5(1'b1), .IN6(na789_1), .IN7(na783_2),
                     .IN8(~na781_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x123y98     80'h00_0018_00_0000_0C66_D500
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1059_1), .IN6(1'b1), .IN7(na2712_2), .IN8(~na2722_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y93     80'h00_0018_00_0000_0666_6C93
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_1 ( .OUT(na791_1), .IN1(1'b0), .IN2(~na2714_2), .IN3(~na1061_1), .IN4(na781_1), .IN5(1'b0), .IN6(na2714_1), .IN7(~na794_1),
                     .IN8(~na1051_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y91     80'h00_0018_00_0040_0AB4_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a794_1 ( .OUT(na794_1), .IN1(1'b1), .IN2(~na2716_2), .IN3(1'b1), .IN4(na781_2), .IN5(na3095_2), .IN6(na2716_1), .IN7(1'b1),
                     .IN8(na1051_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x121y95     80'h00_0060_00_0000_0C08_FF39
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a795_4 ( .OUT(na795_2), .IN1(~na1059_1), .IN2(~na1063_1), .IN3(1'b0), .IN4(na3094_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x121y102     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_1 ( .OUT(na796_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na781_1), .IN5(~na1055_1), .IN6(1'b0), .IN7(~na1053_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y103     80'h00_0018_00_0040_0AF2_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1), .IN1(1'b1), .IN2(~na3197_2), .IN3(~na3099_2), .IN4(1'b1), .IN5(na2718_1), .IN6(~na3164_2), .IN7(na791_1),
                     .IN8(na1461_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y95     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a800_1 ( .OUT(na800_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1055_1), .IN6(na1057_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y106     80'h00_0018_00_0040_0ABD_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a801_1 ( .OUT(na801_1), .IN1(1'b1), .IN2(na802_1), .IN3(1'b1), .IN4(na3103_2), .IN5(~na804_1), .IN6(na2719_2), .IN7(1'b1),
                     .IN8(~na806_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y96     80'h00_0018_00_0040_0AF4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a802_1 ( .OUT(na802_1), .IN1(1'b1), .IN2(~na3164_2), .IN3(~na791_1), .IN4(1'b1), .IN5(na786_1), .IN6(na3197_2), .IN7(~na3198_2),
                     .IN8(na2720_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y99     80'h00_0018_00_0040_0AFA_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a803_1 ( .OUT(na803_1), .IN1(~na786_1), .IN2(1'b1), .IN3(~na791_1), .IN4(1'b1), .IN5(na2718_2), .IN6(~na3197_2), .IN7(na2721_2),
                     .IN8(~na1461_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y105     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a804_1 ( .OUT(na804_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na2729_2), .IN8(na1051_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y108     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a806_1 ( .OUT(na806_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1055_1), .IN6(1'b0), .IN7(~na1053_1), .IN8(na781_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y96     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a807_4 ( .OUT(na807_2), .IN1(~na811_1), .IN2(na809_1), .IN3(~na810_1), .IN4(na808_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y88     80'h00_0018_00_0040_0AE5_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a808_1 ( .OUT(na808_1), .IN1(~na778_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2722_2), .IN5(1'b1), .IN6(na2716_2), .IN7(~na3102_2),
                     .IN8(na2722_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y92     80'h00_0018_00_0040_0AE7_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(~na803_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na781_2), .IN5(1'b1), .IN6(~na3096_2), .IN7(~na797_1),
                     .IN8(na2723_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y103     80'h00_0018_00_0040_0A71_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a810_1 ( .OUT(na810_1), .IN1(1'b1), .IN2(~na3096_2), .IN3(1'b1), .IN4(na781_2), .IN5(~na778_1), .IN6(na2724_1), .IN7(na797_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y91     80'h00_0018_00_0040_0A7E_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a811_1 ( .OUT(na811_1), .IN1(1'b1), .IN2(~na802_1), .IN3(1'b1), .IN4(na3103_2), .IN5(na2725_2), .IN6(~na3101_2), .IN7(~na812_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y87     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a812_1 ( .OUT(na812_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2716_2), .IN7(1'b0), .IN8(na2722_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x121y91     80'h00_0018_00_0000_0C66_7EFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a814_1 ( .OUT(na814_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na803_1), .IN6(~na3097_2), .IN7(na3102_2),
                     .IN8(na781_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y90     80'h00_0018_00_0040_0AB5_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a815_1 ( .OUT(na815_1), .IN1(~na778_1), .IN2(1'b1), .IN3(~na797_1), .IN4(1'b1), .IN5(~na3106_2), .IN6(na2716_2), .IN7(1'b1),
                     .IN8(na2722_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x124y87     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a816_4 ( .OUT(na816_2), .IN1(na818_1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y92     80'h00_0018_00_0040_0A7E_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1), .IN1(na778_1), .IN2(1'b1), .IN3(na2729_2), .IN4(1'b1), .IN5(na3199_2), .IN6(~na802_1), .IN7(~na3142_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y103     80'h00_0018_00_0040_0AE7_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a818_1 ( .OUT(na818_1), .IN1(~na803_1), .IN2(1'b1), .IN3(na797_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2724_2), .IN7(~na3104_2),
                     .IN8(na2730_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x103y98     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a819_1 ( .OUT(na819_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b0), .IN6(na774_1), .IN7(1'b0), .IN8(na2731_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a819_2 ( .OUT(na819_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na819_1_i) );
// C_XOR////D      x113y98     80'h40_E818_00_0000_0666_C590
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a820_1 ( .OUT(na820_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na824_1), .IN4(na776_2), .IN5(~na827_1), .IN6(1'b0), .IN7(1'b0), .IN8(na821_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a820_5 ( .OUT(na820_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na820_1) );
// C_XOR////      x120y100     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a821_1 ( .OUT(na821_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na822_1), .IN6(na809_1), .IN7(na3107_2), .IN8(na808_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y103     80'h00_0018_00_0040_0AB2_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a822_1 ( .OUT(na822_1), .IN1(~na803_1), .IN2(1'b1), .IN3(~na797_1), .IN4(1'b1), .IN5(na804_1), .IN6(~na2719_2), .IN7(1'b0),
                     .IN8(na806_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y104     80'h00_0018_00_0040_0A7A_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a823_1 ( .OUT(na823_1), .IN1(na778_1), .IN2(1'b1), .IN3(~na3102_2), .IN4(1'b1), .IN5(na2733_1), .IN6(~na2724_2), .IN7(na2729_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y101     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a824_1 ( .OUT(na824_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na814_1), .IN6(na815_1), .IN7(~na826_1), .IN8(~na825_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y108     80'h00_0018_00_0040_0AD3_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a825_1 ( .OUT(na825_1), .IN1(1'b1), .IN2(~na802_1), .IN3(1'b1), .IN4(~na3103_2), .IN5(~na804_1), .IN6(1'b1), .IN7(na2734_2),
                     .IN8(na2706_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y107     80'h00_0018_00_0040_0A7E_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a826_1 ( .OUT(na826_1), .IN1(1'b1), .IN2(~na2724_2), .IN3(1'b1), .IN4(~na806_1), .IN5(na778_1), .IN6(~na2724_1), .IN7(~na797_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y99     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na818_1), .IN6(na817_1), .IN7(~na810_1), .IN8(~na3105_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x113y92     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a828_1 ( .OUT(na828_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b0), .IN6(na820_1), .IN7(1'b0), .IN8(na2736_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a828_2 ( .OUT(na828_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na828_1_i) );
// C_XOR////D      x93y109     80'h40_E818_00_0000_0666_0C05
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a829_1 ( .OUT(na829_1), .IN1(~na830_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na831_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a829_5 ( .OUT(na829_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na829_1) );
// C_///XOR/      x113y107     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a830_4 ( .OUT(na830_2), .IN1(na3091_2), .IN2(1'b0), .IN3(na824_1), .IN4(na821_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x111y104     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a831_1 ( .OUT(na831_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na827_1), .IN6(1'b0), .IN7(na824_1), .IN8(na776_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x93y110     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a832_1 ( .OUT(na832_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na829_1), .IN6(1'b0), .IN7(na2737_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a832_2 ( .OUT(na832_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na832_1_i) );
// C_XOR////D      x97y108     80'h40_E818_00_0000_0666_0A30
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a833_1 ( .OUT(na833_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(~na775_1), .IN5(na834_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a833_5 ( .OUT(na833_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na833_1) );
// C_///XOR/      x115y107     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a834_4 ( .OUT(na834_2), .IN1(~na827_1), .IN2(na3108_2), .IN3(na837_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y93     80'h00_0018_00_0040_0ABD_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a836_1 ( .OUT(na836_1), .IN1(~na778_1), .IN2(1'b1), .IN3(~na797_1), .IN4(1'b1), .IN5(~na800_1), .IN6(na2738_1), .IN7(1'b1),
                     .IN8(~na781_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y91     80'h00_0018_00_0040_0AB5_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a837_1 ( .OUT(na837_1), .IN1(1'b1), .IN2(na802_1), .IN3(1'b1), .IN4(na3103_2), .IN5(~na3106_2), .IN6(na2739_2), .IN7(1'b1),
                     .IN8(na781_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x97y99     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a838_1 ( .OUT(na838_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b0), .IN6(na833_1), .IN7(1'b0), .IN8(na2740_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a838_2 ( .OUT(na838_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na838_1_i) );
// C_XOR////D      x101y109     80'h40_E818_00_0000_0666_C005
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_1 ( .OUT(na839_1), .IN1(~na834_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na840_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a839_5 ( .OUT(na839_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na839_1) );
// C_XOR////      x116y102     80'h00_0018_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a840_1 ( .OUT(na840_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na822_1), .IN6(~na823_1), .IN7(na824_1), .IN8(na807_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x100y104     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a841_1 ( .OUT(na841_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na839_1), .IN6(1'b0), .IN7(na2741_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a841_2 ( .OUT(na841_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na841_1_i) );
// C_XOR////D      x117y97     80'h40_E818_00_0000_0666_999A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a842_1 ( .OUT(na842_1), .IN1(na822_1), .IN2(1'b0), .IN3(~na824_1), .IN4(na776_2), .IN5(~na836_1), .IN6(na823_1), .IN7(~na837_1),
                     .IN8(na807_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a842_5 ( .OUT(na842_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na842_1) );
// C_MX2b/D///      x104y89     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a844_1 ( .OUT(na844_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na842_1), .IN6(1'b0), .IN7(na2742_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a844_2 ( .OUT(na844_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na844_1_i) );
// C_XOR////D      x120y91     80'h40_E818_00_0000_0666_0996
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a845_1 ( .OUT(na845_1), .IN1(na836_1), .IN2(na815_1), .IN3(na837_1), .IN4(~na808_1), .IN5(na814_1), .IN6(~na809_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a845_5 ( .OUT(na845_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na845_1) );
// C_MX2b/D///      x107y88     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a846_1 ( .OUT(na846_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na2743_2), .IN6(1'b0), .IN7(na845_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a846_2 ( .OUT(na846_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na846_1_i) );
// C_XOR////D      x117y101     80'h40_E818_00_0000_0666_999A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_1 ( .OUT(na847_1), .IN1(na822_1), .IN2(1'b0), .IN3(~na824_1), .IN4(na776_2), .IN5(~na836_1), .IN6(na823_1), .IN7(~na837_1),
                     .IN8(na821_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a847_5 ( .OUT(na847_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na847_1) );
// C_MX2b/D///      x99y102     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a848_1 ( .OUT(na848_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na847_1), .IN6(1'b0), .IN7(na2744_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a848_2 ( .OUT(na848_1), .CLK(1'b0), .EN(na1109_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na848_1_i) );
// C_XOR////D      x87y103     80'h40_E818_00_0000_0666_0CA0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a849_1 ( .OUT(na849_1), .IN1(1'b0), .IN2(1'b0), .IN3(na850_1), .IN4(1'b0), .IN5(1'b0), .IN6(na895_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a849_5 ( .OUT(na849_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na849_1) );
// C_XOR////      x110y109     80'h00_0018_00_0000_0666_A9AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a850_1 ( .OUT(na850_1), .IN1(1'b0), .IN2(na2766_2), .IN3(na851_1), .IN4(1'b0), .IN5(na894_1), .IN6(~na2766_1), .IN7(na851_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x116y101     80'h00_0078_00_0000_0C66_AC96
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a851_1 ( .OUT(na851_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na852_1), .IN7(na881_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a851_4 ( .OUT(na851_2), .IN1(na891_1), .IN2(na888_1), .IN3(na889_1), .IN4(~na890_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y110     80'h00_0018_00_0040_0A76_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a852_1 ( .OUT(na852_1), .IN1(na853_1), .IN2(1'b1), .IN3(na877_1), .IN4(1'b1), .IN5(na2745_2), .IN6(~na879_2), .IN7(~na878_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y109     80'h00_0018_00_0040_0AF2_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_1 ( .OUT(na853_1), .IN1(na1465_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3118_2), .IN5(na2746_1), .IN6(~na3200_2), .IN7(na2758_2),
                     .IN8(na868_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x115y107     80'h00_0018_00_0000_0C66_6300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a856_1 ( .OUT(na856_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1079_1), .IN7(na3146_2), .IN8(na1075_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x116y110     80'h00_0078_00_0000_0C66_A569
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a858_1 ( .OUT(na858_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1071_1), .IN6(1'b0), .IN7(na1069_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a858_4 ( .OUT(na858_2), .IN1(na3148_2), .IN2(~na1079_1), .IN3(na1069_1), .IN4(na1075_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x115y110     80'h00_0078_00_0000_0C66_99C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a860_1 ( .OUT(na860_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1071_1), .IN6(~na1077_1), .IN7(na1073_1),
                     .IN8(~na1081_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a860_4 ( .OUT(na860_2), .IN1(1'b0), .IN2(~na1077_1), .IN3(1'b0), .IN4(na1081_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y104     80'h00_0018_00_0040_0A98_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a862_1 ( .OUT(na862_1), .IN1(na1071_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3147_2), .IN5(na3148_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na1081_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x121y108     80'h00_0018_00_0000_0666_3D57
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a863_1 ( .OUT(na863_1), .IN1(na2750_1), .IN2(na860_1), .IN3(na865_1), .IN4(1'b1), .IN5(na2750_2), .IN6(~na860_2), .IN7(1'b1),
                     .IN8(na1075_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x116y109     80'h00_0018_00_0040_0AD9_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a865_1 ( .OUT(na865_1), .IN1(na3201_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na858_2), .IN5(~na856_1), .IN6(1'b0), .IN7(na2751_1),
                     .IN8(~na858_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x118y110     80'h00_0018_00_0000_0666_EE57
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_1 ( .OUT(na868_1), .IN1(na3201_2), .IN2(na860_1), .IN3(na869_1), .IN4(1'b1), .IN5(~na3112_2), .IN6(~na860_2), .IN7(~na2757_2),
                     .IN8(~na858_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y105     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1), .IN1(1'b1), .IN2(na1067_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na870_2), .IN6(~na1077_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x117y103     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a870_4 ( .OUT(na870_2), .IN1(1'b0), .IN2(na1079_1), .IN3(1'b0), .IN4(~na1075_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x118y109     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a874_1 ( .OUT(na874_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3116_2), .IN5(na2756_2), .IN6(1'b0), .IN7(na2757_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y109     80'h00_0018_00_0040_0AB2_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_1 ( .OUT(na875_1), .IN1(1'b1), .IN2(~na3203_2), .IN3(na2751_2), .IN4(1'b1), .IN5(na870_2), .IN6(~na1077_1), .IN7(1'b0),
                     .IN8(na3202_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y110     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a876_1 ( .OUT(na876_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na3115_2), .IN5(~na1071_1), .IN6(1'b0), .IN7(~na1069_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y109     80'h00_0018_00_0040_0AF2_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_1 ( .OUT(na877_1), .IN1(1'b1), .IN2(~na863_1), .IN3(na2758_2), .IN4(1'b1), .IN5(na1465_1), .IN6(~na3165_2), .IN7(na2758_1),
                     .IN8(na868_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x122y105     80'h00_0078_00_0000_0C66_06CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_1 ( .OUT(na878_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3201_2), .IN6(na860_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a878_4 ( .OUT(na878_2), .IN1(1'b0), .IN2(na3113_2), .IN3(1'b0), .IN4(na858_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y110     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a879_4 ( .OUT(na879_2), .IN1(~na2750_2), .IN2(1'b0), .IN3(1'b0), .IN4(na880_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x112y108     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a880_1 ( .OUT(na880_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1071_1), .IN6(1'b0), .IN7(na1073_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y109     80'h00_0018_00_0040_0A7E_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a881_1 ( .OUT(na881_1), .IN1(1'b1), .IN2(~na3123_2), .IN3(1'b1), .IN4(na3124_2), .IN5(na2759_1), .IN6(~na3125_2), .IN7(~na878_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y108     80'h00_0018_00_0040_0AF4_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a882_1 ( .OUT(na882_1), .IN1(~na1465_1), .IN2(1'b1), .IN3(1'b1), .IN4(na868_1), .IN5(na3117_2), .IN6(na3204_2), .IN7(~na2758_2),
                     .IN8(na2760_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y108     80'h00_0018_00_0040_0AF5_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_1 ( .OUT(na883_1), .IN1(1'b1), .IN2(na3204_2), .IN3(1'b1), .IN4(na868_1), .IN5(~na3117_2), .IN6(na863_1), .IN7(~na3166_2),
                     .IN8(na2761_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y105     80'h00_0018_00_0000_0C66_5C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a884_1 ( .OUT(na884_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1067_1), .IN7(~na2769_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y106     80'h00_0018_00_0040_0ADA_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a888_1 ( .OUT(na888_1), .IN1(na853_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3116_2), .IN5(na856_1), .IN6(1'b1), .IN7(na2762_2),
                     .IN8(~na882_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y103     80'h00_0018_00_0040_0AE3_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a889_1 ( .OUT(na889_1), .IN1(1'b1), .IN2(~na883_1), .IN3(~na877_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na860_1), .IN7(na3114_2),
                     .IN8(na3205_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y110     80'h00_0018_00_0040_0AB9_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a890_1 ( .OUT(na890_1), .IN1(~na853_1), .IN2(1'b1), .IN3(na877_1), .IN4(1'b1), .IN5(~na2763_1), .IN6(na860_1), .IN7(1'b0),
                     .IN8(~na858_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y107     80'h00_0018_00_0040_0ABD_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1), .IN1(1'b1), .IN2(~na883_1), .IN3(1'b1), .IN4(~na882_1), .IN5(~na892_1), .IN6(na2765_2), .IN7(1'b1),
                     .IN8(~na880_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y107     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a892_1 ( .OUT(na892_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na856_1), .IN6(na860_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x115y105     80'h00_0018_00_0040_0A7C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a894_1 ( .OUT(na894_1), .IN1(na3119_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3111_2), .IN5(na856_1), .IN6(na860_2), .IN7(~na3126_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x107y110     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a895_4 ( .OUT(na895_2), .IN1(na896_1), .IN2(1'b0), .IN3(na897_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y109     80'h00_0018_00_0040_0ADB_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a896_1 ( .OUT(na896_1), .IN1(na853_1), .IN2(1'b1), .IN3(~na2769_2), .IN4(1'b1), .IN5(~na3145_2), .IN6(1'b1), .IN7(na2769_1),
                     .IN8(~na882_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y107     80'h00_0018_00_0040_0AE5_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1), .IN1(1'b1), .IN2(~na883_1), .IN3(~na877_1), .IN4(1'b1), .IN5(1'b1), .IN6(na3120_2), .IN7(~na878_2),
                     .IN8(na2770_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x91y98     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a898_1 ( .OUT(na898_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na849_1), .IN6(1'b0), .IN7(na2771_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a898_2 ( .OUT(na898_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na898_1_i) );
// C_XOR////D      x98y110     80'h40_E818_00_0000_0666_390A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a899_1 ( .OUT(na899_1), .IN1(na900_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na891_1), .IN6(na895_2), .IN7(1'b0), .IN8(~na890_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a899_5 ( .OUT(na899_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na899_1) );
// C_XOR///XOR/      x111y101     80'h00_0078_00_0000_0C66_6960
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_1 ( .OUT(na900_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1467_1), .IN6(na904_1), .IN7(na851_1), .IN8(na901_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a900_4 ( .OUT(na900_2), .IN1(1'b0), .IN2(1'b0), .IN3(na906_1), .IN4(na3127_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x110y108     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a901_1 ( .OUT(na901_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na888_1), .IN7(na889_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y102     80'h00_0018_00_0000_0666_A65C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a904_1 ( .OUT(na904_1), .IN1(1'b0), .IN2(na2766_2), .IN3(~na905_1), .IN4(1'b0), .IN5(na894_1), .IN6(na2766_1), .IN7(na906_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y101     80'h00_0018_00_0040_0ADC_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a905_1 ( .OUT(na905_1), .IN1(na853_1), .IN2(1'b1), .IN3(~na877_1), .IN4(1'b1), .IN5(na3121_2), .IN6(1'b0), .IN7(~na878_1),
                     .IN8(~na2770_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y103     80'h00_0018_00_0040_0AE5_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a906_1 ( .OUT(na906_1), .IN1(1'b1), .IN2(~na883_1), .IN3(1'b1), .IN4(na882_1), .IN5(1'b1), .IN6(na879_2), .IN7(~na884_1),
                     .IN8(na2773_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x98y107     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a907_1 ( .OUT(na907_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na429_1), .IN5(1'b0), .IN6(na2774_2), .IN7(1'b0), .IN8(na899_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a907_2 ( .OUT(na907_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na907_1_i) );
// C_XOR////D      x99y110     80'h40_E818_00_0000_0666_CAA6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a908_1 ( .OUT(na908_1), .IN1(~na900_2), .IN2(~na895_2), .IN3(na850_1), .IN4(1'b0), .IN5(na900_1), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na901_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a908_5 ( .OUT(na908_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na908_1) );
// C_MX2b/D///      x95y103     80'h40_E800_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a911_1 ( .OUT(na911_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b0), .IN6(na908_1), .IN7(1'b0), .IN8(na3208_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a911_2 ( .OUT(na911_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na911_1_i) );
// C_XOR////D      x98y97     80'h40_E818_00_0000_0666_A030
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a912_1 ( .OUT(na912_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(~na913_1), .IN5(1'b0), .IN6(1'b0), .IN7(na850_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a912_5 ( .OUT(na912_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na912_1) );
// C_XOR////      x114y102     80'h00_0018_00_0000_0666_9666
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a913_1 ( .OUT(na913_1), .IN1(na3110_2), .IN2(na895_2), .IN3(na905_1), .IN4(na901_1), .IN5(~na900_2), .IN6(~na916_1), .IN7(na906_1),
                     .IN8(~na915_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y104     80'h00_0018_00_0040_0AD8_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a915_1 ( .OUT(na915_1), .IN1(1'b1), .IN2(na883_1), .IN3(1'b1), .IN4(na882_1), .IN5(na892_1), .IN6(1'b0), .IN7(na2776_2),
                     .IN8(~na858_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y104     80'h00_0018_00_0040_0AE7_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a916_1 ( .OUT(na916_1), .IN1(~na853_1), .IN2(1'b1), .IN3(~na877_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na860_1), .IN7(~na3122_2),
                     .IN8(na2777_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x94y92     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a917_1 ( .OUT(na917_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na2778_2), .IN6(1'b0), .IN7(na912_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a917_2 ( .OUT(na917_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na917_1_i) );
// C_XOR////D      x102y99     80'h40_E818_00_0000_0666_A030
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a918_1 ( .OUT(na918_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(~na913_1), .IN5(1'b0), .IN6(1'b0), .IN7(na919_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a918_5 ( .OUT(na918_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na918_1) );
// C_///XOR/      x118y101     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a919_4 ( .OUT(na919_2), .IN1(na1467_1), .IN2(~na904_1), .IN3(na851_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x100y92     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_1 ( .OUT(na920_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na2779_1), .IN6(1'b0), .IN7(na918_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a920_2 ( .OUT(na920_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na920_1_i) );
// C_XOR////D      x117y85     80'h40_E818_00_0000_0666_605A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a921_1 ( .OUT(na921_1), .IN1(na900_2), .IN2(1'b0), .IN3(~na851_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na851_2), .IN8(na923_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a921_5 ( .OUT(na921_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na921_1) );
// C_XOR////      x114y100     80'h00_0018_00_0000_0666_AC99
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a923_1 ( .OUT(na923_1), .IN1(na1467_1), .IN2(~na916_1), .IN3(na905_1), .IN4(~na915_1), .IN5(1'b0), .IN6(na904_1), .IN7(na906_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x104y84     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a924_1 ( .OUT(na924_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na921_1), .IN6(1'b0), .IN7(na2780_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a924_2 ( .OUT(na924_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na924_1_i) );
// C_XOR////D      x103y73     80'h40_E818_00_0000_0666_CAC0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a925_1 ( .OUT(na925_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na923_1), .IN5(na1467_1), .IN6(1'b0), .IN7(1'b0), .IN8(na901_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a925_5 ( .OUT(na925_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na925_1) );
// C_MX2b/D///      x99y76     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a926_1 ( .OUT(na926_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na925_1), .IN6(1'b0), .IN7(na2781_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a926_2 ( .OUT(na926_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na926_1_i) );
// C_XOR////D      x109y81     80'h40_E818_00_0000_0666_9AA5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a927_1 ( .OUT(na927_1), .IN1(~na900_1), .IN2(1'b0), .IN3(na851_2), .IN4(1'b0), .IN5(na3109_2), .IN6(1'b0), .IN7(~na851_1),
                     .IN8(na923_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a927_5 ( .OUT(na927_2), .CLK(1'b0), .EN(na1108_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na927_1) );
// C_MX2b/D///      x102y82     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a928_1 ( .OUT(na928_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na927_1), .IN6(1'b0), .IN7(na2782_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a928_2 ( .OUT(na928_1), .CLK(1'b0), .EN(na1110_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na928_1_i) );
// C_MX2b/D///      x110y87     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a929_1 ( .OUT(na929_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na2691_1), .IN6(1'b0), .IN7(na693_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a929_2 ( .OUT(na929_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na929_1_i) );
// C_MX2b/D///      x104y94     80'h40_E800_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a930_1 ( .OUT(na930_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na739_1), .IN6(1'b0), .IN7(na2697_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a930_2 ( .OUT(na930_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na930_1_i) );
// C_MX2b/D///      x104y88     80'h40_E800_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a931_1 ( .OUT(na931_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na748_1), .IN6(1'b0), .IN7(na2698_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a931_2 ( .OUT(na931_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na931_1_i) );
// C_MX2b/D///      x101y80     80'h40_E800_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a932_1 ( .OUT(na932_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na754_1), .IN6(1'b0), .IN7(na2701_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a932_2 ( .OUT(na932_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na932_1_i) );
// C_MX2b/D///      x100y80     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a933_1 ( .OUT(na933_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na2702_2), .IN6(1'b0), .IN7(na760_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a933_2 ( .OUT(na933_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na933_1_i) );
// C_MX2b/D///      x103y69     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a934_1 ( .OUT(na934_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na2703_1), .IN6(1'b0), .IN7(na764_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a934_2 ( .OUT(na934_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na934_1_i) );
// C_MX2b/D///      x102y74     80'h40_E800_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a935_1 ( .OUT(na935_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na769_1), .IN6(1'b0), .IN7(na2704_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a935_2 ( .OUT(na935_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na935_1_i) );
// C_MX2b/D///      x101y74     80'h40_E800_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a936_1 ( .OUT(na936_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na771_1), .IN7(1'b0), .IN8(na3195_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a936_2 ( .OUT(na936_1), .CLK(1'b0), .EN(na1105_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na936_1_i) );
// C_MX2b/D///      x102y98     80'h40_E400_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a937_1 ( .OUT(na937_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na774_1), .IN7(1'b0), .IN8(na2731_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a937_2 ( .OUT(na937_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na937_1_i) );
// C_MX2b/D///      x106y94     80'h40_E400_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a938_1 ( .OUT(na938_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na820_1), .IN7(1'b0), .IN8(na2736_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a938_2 ( .OUT(na938_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na938_1_i) );
// C_MX2b/D///      x91y107     80'h40_E400_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a939_1 ( .OUT(na939_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na829_1), .IN6(1'b0), .IN7(na2737_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a939_2 ( .OUT(na939_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na939_1_i) );
// C_MX2b/D///      x96y104     80'h40_E400_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a940_1 ( .OUT(na940_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na833_1), .IN7(1'b0), .IN8(na2740_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a940_2 ( .OUT(na940_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na940_1_i) );
// C_MX2b/D///      x99y100     80'h40_E400_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a941_1 ( .OUT(na941_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na839_1), .IN6(1'b0), .IN7(na2741_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a941_2 ( .OUT(na941_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na941_1_i) );
// C_MX2b/D///      x110y92     80'h40_E400_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a942_1 ( .OUT(na942_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na842_1), .IN6(1'b0), .IN7(na2742_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a942_2 ( .OUT(na942_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na942_1_i) );
// C_MX2b/D///      x113y87     80'h40_E400_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a943_1 ( .OUT(na943_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na2743_2), .IN6(1'b0), .IN7(na845_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a943_2 ( .OUT(na943_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na943_1_i) );
// C_MX2b/D///      x103y102     80'h40_E400_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a944_1 ( .OUT(na944_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na847_1), .IN6(1'b0), .IN7(na2744_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a944_2 ( .OUT(na944_1), .CLK(1'b0), .EN(~na1100_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na944_1_i) );
// C_MX2b/D///      x91y97     80'h40_E400_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_1 ( .OUT(na945_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na849_1), .IN6(1'b0), .IN7(na2771_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a945_2 ( .OUT(na945_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na945_1_i) );
// C_MX2b/D///      x93y106     80'h40_E400_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a946_1 ( .OUT(na946_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b0), .IN6(na2774_2), .IN7(1'b0), .IN8(na899_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a946_2 ( .OUT(na946_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na946_1_i) );
// C_MX2b/D///      x94y103     80'h40_E400_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a947_1 ( .OUT(na947_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na429_1), .IN5(1'b0), .IN6(na908_1), .IN7(1'b0), .IN8(na3208_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a947_2 ( .OUT(na947_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na947_1_i) );
// C_MX2b/D///      x95y92     80'h40_E400_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a948_1 ( .OUT(na948_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na2778_2), .IN6(1'b0), .IN7(na912_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a948_2 ( .OUT(na948_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na948_1_i) );
// C_MX2b/D///      x99y90     80'h40_E400_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a949_1 ( .OUT(na949_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na2779_1), .IN6(1'b0), .IN7(na918_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a949_2 ( .OUT(na949_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na949_1_i) );
// C_MX2b/D///      x103y84     80'h40_E400_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a950_1 ( .OUT(na950_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na921_1), .IN6(1'b0), .IN7(na2780_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a950_2 ( .OUT(na950_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na950_1_i) );
// C_MX2b/D///      x99y74     80'h40_E400_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a951_1 ( .OUT(na951_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na925_1), .IN6(1'b0), .IN7(na2781_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a951_2 ( .OUT(na951_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na951_1_i) );
// C_MX2b/D///      x99y84     80'h40_E400_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a952_1 ( .OUT(na952_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na927_1), .IN6(1'b0), .IN7(na2782_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a952_2 ( .OUT(na952_1), .CLK(1'b0), .EN(~na1095_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na952_1_i) );
// C_MX2b/D///      x112y82     80'h40_E400_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a953_1 ( .OUT(na953_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na693_1), .IN8(na3185_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a953_2 ( .OUT(na953_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na953_1_i) );
// C_MX2b/D///      x105y91     80'h40_E400_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a954_1 ( .OUT(na954_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na739_1), .IN6(na3189_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a954_2 ( .OUT(na954_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na954_1_i) );
// C_MX2b/D///      x107y82     80'h40_E400_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a955_1 ( .OUT(na955_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na748_1), .IN6(na3190_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a955_2 ( .OUT(na955_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na955_1_i) );
// C_MX2b/D///      x101y78     80'h40_E400_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a956_1 ( .OUT(na956_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na754_1), .IN6(na3191_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a956_2 ( .OUT(na956_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na956_1_i) );
// C_MX2b/D///      x101y77     80'h40_E400_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a957_1 ( .OUT(na957_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na760_1), .IN8(na3192_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a957_2 ( .OUT(na957_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na957_1_i) );
// C_MX2b/D///      x107y69     80'h40_E400_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a958_1 ( .OUT(na958_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na764_1), .IN8(na3193_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a958_2 ( .OUT(na958_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na958_1_i) );
// C_MX2b/D///      x101y70     80'h40_E400_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a959_1 ( .OUT(na959_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na769_1), .IN6(na3194_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a959_2 ( .OUT(na959_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na959_1_i) );
// C_MX2b/D///      x103y71     80'h40_E400_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a960_1 ( .OUT(na960_1_i), .IN1(1'b1), .IN2(~na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2705_1), .IN6(na771_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a960_2 ( .OUT(na960_1), .CLK(1'b0), .EN(~na1098_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na960_1_i) );
// C_MX2b/D///      x105y96     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a961_1 ( .OUT(na961_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na429_1), .IN5(1'b0), .IN6(na774_1), .IN7(1'b0), .IN8(na2731_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a961_2 ( .OUT(na961_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na961_1_i) );
// C_MX2b/D///      x109y91     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a962_1 ( .OUT(na962_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na429_1), .IN5(1'b0), .IN6(na820_1), .IN7(1'b0), .IN8(na2736_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a962_2 ( .OUT(na962_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na962_1_i) );
// C_MX2b/D///      x91y104     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a963_1 ( .OUT(na963_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na829_1), .IN6(1'b0), .IN7(na2737_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a963_2 ( .OUT(na963_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na963_1_i) );
// C_MX2b/D///      x102y102     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a964_1 ( .OUT(na964_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na429_1), .IN5(1'b0), .IN6(na833_1), .IN7(1'b0), .IN8(na2740_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a964_2 ( .OUT(na964_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na964_1_i) );
// C_MX2b/D///      x98y102     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a965_1 ( .OUT(na965_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na839_1), .IN6(1'b0), .IN7(na2741_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a965_2 ( .OUT(na965_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na965_1_i) );
// C_MX2b/D///      x115y90     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a966_1 ( .OUT(na966_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na842_1), .IN6(1'b0), .IN7(na2742_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a966_2 ( .OUT(na966_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na966_1_i) );
// C_MX2b/D///      x113y86     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a967_1 ( .OUT(na967_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na2743_2), .IN6(1'b0), .IN7(na845_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a967_2 ( .OUT(na967_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na967_1_i) );
// C_MX2b/D///      x105y100     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a968_1 ( .OUT(na968_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na847_1), .IN6(1'b0), .IN7(na2744_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a968_2 ( .OUT(na968_1), .CLK(1'b0), .EN(na1094_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na968_1_i) );
// C_MX2b/D///      x93y97     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a969_1 ( .OUT(na969_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na849_1), .IN6(1'b0), .IN7(na2771_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a969_2 ( .OUT(na969_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na969_1_i) );
// C_MX2b/D///      x96y107     80'h40_E800_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a970_1 ( .OUT(na970_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na2774_2), .IN7(1'b0), .IN8(na899_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a970_2 ( .OUT(na970_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na970_1_i) );
// C_MX2b/D///      x95y104     80'h40_E800_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a971_1 ( .OUT(na971_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na908_1), .IN7(1'b0), .IN8(na3208_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a971_2 ( .OUT(na971_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na971_1_i) );
// C_MX2b/D///      x97y95     80'h40_E800_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a972_1 ( .OUT(na972_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na2778_2), .IN6(1'b0), .IN7(na912_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a972_2 ( .OUT(na972_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na972_1_i) );
// C_MX2b/D///      x100y94     80'h40_E800_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_1 ( .OUT(na973_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na2779_1), .IN6(1'b0), .IN7(na918_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a973_2 ( .OUT(na973_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na973_1_i) );
// C_MX2b/D///      x103y86     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a974_1 ( .OUT(na974_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na921_1), .IN6(1'b0), .IN7(na2780_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a974_2 ( .OUT(na974_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na974_1_i) );
// C_MX2b/D///      x100y79     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a975_1 ( .OUT(na975_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na925_1), .IN6(1'b0), .IN7(na2781_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a975_2 ( .OUT(na975_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na975_1_i) );
// C_MX2b/D///      x101y87     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a976_1 ( .OUT(na976_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na927_1), .IN6(1'b0), .IN7(na2782_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a976_2 ( .OUT(na976_1), .CLK(1'b0), .EN(na1106_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na976_1_i) );
// C_MX2b/D///      x111y81     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a977_1 ( .OUT(na977_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na2691_1), .IN6(1'b0), .IN7(na693_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a977_2 ( .OUT(na977_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na977_1_i) );
// C_MX2b/D///      x105y90     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a978_1 ( .OUT(na978_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na739_1), .IN6(1'b0), .IN7(na2697_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a978_2 ( .OUT(na978_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na978_1_i) );
// C_MX2b/D///      x109y84     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a979_1 ( .OUT(na979_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na748_1), .IN6(1'b0), .IN7(na2698_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a979_2 ( .OUT(na979_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na979_1_i) );
// C_MX2b/D///      x107y80     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a980_1 ( .OUT(na980_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na754_1), .IN6(1'b0), .IN7(na2701_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a980_2 ( .OUT(na980_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na980_1_i) );
// C_MX2b/D///      x102y78     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a981_1 ( .OUT(na981_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na2702_2), .IN6(1'b0), .IN7(na760_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a981_2 ( .OUT(na981_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na981_1_i) );
// C_MX2b/D///      x103y66     80'h40_E800_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a982_1 ( .OUT(na982_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_1), .IN5(na2703_1), .IN6(1'b0), .IN7(na764_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a982_2 ( .OUT(na982_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na982_1_i) );
// C_MX2b/D///      x103y70     80'h40_E800_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a983_1 ( .OUT(na983_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na769_1), .IN6(1'b0), .IN7(na2704_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a983_2 ( .OUT(na983_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na983_1_i) );
// C_MX2b/D///      x104y72     80'h40_E800_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a984_1 ( .OUT(na984_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na429_1), .IN5(1'b0), .IN6(na771_1), .IN7(1'b0), .IN8(na3195_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a984_2 ( .OUT(na984_1), .CLK(1'b0), .EN(na1091_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na984_1_i) );
// C_MX2b/D///      x101y98     80'h40_E800_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a985_1 ( .OUT(na985_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na774_1), .IN7(1'b0), .IN8(na2731_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a985_2 ( .OUT(na985_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na985_1_i) );
// C_MX2b/D///      x106y92     80'h40_E800_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a986_1 ( .OUT(na986_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na820_1), .IN7(1'b0), .IN8(na2736_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a986_2 ( .OUT(na986_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na986_1_i) );
// C_MX2b/D///      x93y105     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a987_1 ( .OUT(na987_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na829_1), .IN6(1'b0), .IN7(na2737_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a987_2 ( .OUT(na987_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na987_1_i) );
// C_MX2b/D///      x97y102     80'h40_E800_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a988_1 ( .OUT(na988_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(1'b0), .IN6(na833_1), .IN7(1'b0), .IN8(na2740_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a988_2 ( .OUT(na988_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na988_1_i) );
// C_MX2b/D///      x99y104     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a989_1 ( .OUT(na989_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na839_1), .IN6(1'b0), .IN7(na2741_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a989_2 ( .OUT(na989_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na989_1_i) );
// C_MX2b/D///      x111y92     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a990_1 ( .OUT(na990_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na842_1), .IN6(1'b0), .IN7(na2742_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a990_2 ( .OUT(na990_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na990_1_i) );
// C_MX2b/D///      x111y88     80'h40_E800_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a991_1 ( .OUT(na991_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1103_2), .IN4(1'b1), .IN5(na2743_2), .IN6(1'b0), .IN7(na845_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a991_2 ( .OUT(na991_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na991_1_i) );
// C_MX2b/D///      x104y102     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a992_1 ( .OUT(na992_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b1), .IN5(na847_1), .IN6(1'b0), .IN7(na2744_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a992_2 ( .OUT(na992_1), .CLK(1'b0), .EN(na1101_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na992_1_i) );
// C_MX2b/D///      x90y97     80'h40_E800_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a993_1 ( .OUT(na993_1_i), .IN1(1'b1), .IN2(~na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na849_1), .IN6(na3206_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a993_2 ( .OUT(na993_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na993_1_i) );
// C_MX2b/D///      x93y107     80'h40_E800_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a994_1 ( .OUT(na994_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3207_2), .IN8(na899_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a994_2 ( .OUT(na994_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na994_1_i) );
// C_MX2b/D///      x89y99     80'h40_E800_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_1 ( .OUT(na995_1_i), .IN1(1'b1), .IN2(na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2775_1), .IN6(na908_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a995_2 ( .OUT(na995_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na995_1_i) );
// C_MX2b/D///      x93y92     80'h40_E800_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a996_1 ( .OUT(na996_1_i), .IN1(1'b1), .IN2(~na104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na912_1), .IN8(na3209_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a996_2 ( .OUT(na996_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na996_1_i) );
// C_MX2b/D///      x95y91     80'h40_E800_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a997_1 ( .OUT(na997_1_i), .IN1(1'b1), .IN2(~na104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na918_1), .IN8(na3210_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a997_2 ( .OUT(na997_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na997_1_i) );
// C_MX2b/D///      x101y83     80'h40_E800_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a998_1 ( .OUT(na998_1_i), .IN1(1'b1), .IN2(~na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na921_1), .IN6(na3211_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a998_2 ( .OUT(na998_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na998_1_i) );
// C_MX2b/D///      x98y76     80'h40_E800_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_1 ( .OUT(na999_1_i), .IN1(1'b1), .IN2(~na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na925_1), .IN6(na3212_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a999_2 ( .OUT(na999_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na999_1_i) );
// C_MX2b/D///      x99y82     80'h40_E800_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1_i), .IN1(1'b1), .IN2(~na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(na927_1), .IN6(na3213_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1000_2 ( .OUT(na1000_1), .CLK(1'b0), .EN(na1102_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1000_1_i) );
// C_MX2b/D///      x90y109     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1001_1 ( .OUT(na1001_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na66_1), .IN4(1'b1), .IN5(na11_1), .IN6(1'b0), .IN7(na3214_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1001_2 ( .OUT(na1001_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1001_1_i) );
// C_MX2b/D///      x85y110     80'h40_E800_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1002_1 ( .OUT(na1002_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na66_1), .IN4(1'b1), .IN5(1'b0), .IN6(na2856_1), .IN7(1'b0), .IN8(na69_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1002_2 ( .OUT(na1002_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1002_1_i) );
// C_MX2b/D///      x89y106     80'h40_E800_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_1 ( .OUT(na1003_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b0), .IN6(na85_1), .IN7(1'b0), .IN8(na2857_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1003_2 ( .OUT(na1003_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1003_1_i) );
// C_MX2b/D///      x89y102     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1004_1 ( .OUT(na1004_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na66_1), .IN4(1'b1), .IN5(na94_1), .IN6(1'b0), .IN7(na2858_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1004_2 ( .OUT(na1004_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1004_1_i) );
// C_MX2b/D///      x90y99     80'h40_E800_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1005_1 ( .OUT(na1005_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b0), .IN6(na105_1), .IN7(1'b0), .IN8(na2859_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1005_2 ( .OUT(na1005_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1005_1_i) );
// C_MX2b/D///      x95y95     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1006_1 ( .OUT(na1006_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na66_1), .IN4(1'b1), .IN5(na112_1), .IN6(1'b0), .IN7(na2860_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1006_2 ( .OUT(na1006_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1006_1_i) );
// C_MX2b/D///      x100y95     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1007_1 ( .OUT(na1007_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na66_1), .IN4(1'b1), .IN5(na121_1), .IN6(1'b0), .IN7(na2861_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1007_2 ( .OUT(na1007_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1007_1_i) );
// C_MX2b/D///      x96y98     80'h40_E800_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1008_1 ( .OUT(na1008_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na66_1), .IN4(1'b1), .IN5(na128_1), .IN6(1'b0), .IN7(na2862_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1008_2 ( .OUT(na1008_1), .CLK(1'b0), .EN(na1107_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1008_1_i) );
// C_MX2b////D      x85y99     80'h40_E818_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1010_1), .IN5(na11_1), .IN6(1'b0), .IN7(na3214_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1009_5 ( .OUT(na1009_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1009_1) );
// C_AND///AND/      x96y88     80'h00_0078_00_0000_0C88_8431
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_1 ( .OUT(na1010_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1087_2), .IN6(na1090_2), .IN7(na1089_2),
                      .IN8(na3158_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1010_4 ( .OUT(na1010_2), .IN1(~na1087_2), .IN2(~na2923_2), .IN3(1'b1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x83y103     80'h40_E818_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1011_1 ( .OUT(na1011_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1010_1), .IN5(1'b0), .IN6(na2856_1), .IN7(1'b0), .IN8(na69_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1011_5 ( .OUT(na1011_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1011_1) );
// C_MX2b////D      x85y93     80'h40_E818_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_1 ( .OUT(na1012_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1010_1), .IN5(1'b0), .IN6(na85_1), .IN7(1'b0), .IN8(na2857_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1012_5 ( .OUT(na1012_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1012_1) );
// C_MX2b////D      x85y84     80'h40_E818_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1013_1 ( .OUT(na1013_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1010_1), .IN5(na94_1), .IN6(1'b0), .IN7(na2858_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1013_5 ( .OUT(na1013_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1013_1) );
// C_MX2b////D      x87y79     80'h40_E818_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1014_1 ( .OUT(na1014_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1010_1), .IN5(1'b0), .IN6(na105_1), .IN7(1'b0), .IN8(na2859_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1014_5 ( .OUT(na1014_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1014_1) );
// C_MX2b////D      x92y71     80'h40_E818_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1015_1 ( .OUT(na1015_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1010_1), .IN5(na112_1), .IN6(1'b0), .IN7(na2860_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1015_5 ( .OUT(na1015_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1015_1) );
// C_MX2b////D      x90y75     80'h40_E818_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_1 ( .OUT(na1016_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1010_1), .IN5(na121_1), .IN6(1'b0), .IN7(na2861_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1016_5 ( .OUT(na1016_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1016_1) );
// C_MX2b////D      x87y75     80'h40_E818_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1017_1 ( .OUT(na1017_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1010_1), .IN5(na128_1), .IN6(1'b0), .IN7(na2862_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1017_5 ( .OUT(na1017_2), .CLK(1'b0), .EN(na65_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1017_1) );
// C_MX2b/D///      x84y91     80'h40_EC00_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_1 ( .OUT(na1018_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1020_1), .IN6(na2855_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1018_2 ( .OUT(na1018_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1018_1_i) );
// C_MX2b////      x89y95     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1020_1 ( .OUT(na1020_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na428_1), .IN8(~na461_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x82y98     80'h40_EC00_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1021_1 ( .OUT(na1021_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1022_1), .IN6(na2856_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1021_2 ( .OUT(na1021_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1021_1_i) );
// C_MX2b////      x85y101     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_1 ( .OUT(na1022_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na430_1), .IN6(~na462_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x81y96     80'h40_EC00_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_1 ( .OUT(na1023_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1024_1),
                      .IN8(na2857_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1023_2 ( .OUT(na1023_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1023_1_i) );
// C_MX2b////      x88y93     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1024_1 ( .OUT(na1024_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na463_2), .IN6(~na431_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x86y89     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2858_1), .IN8(~na1026_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1025_2 ( .OUT(na1025_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1025_1_i) );
// C_MX2b////      x92y84     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1026_1 ( .OUT(na1026_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na432_2), .IN6(~na464_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x82y93     80'h40_EC00_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1027_1 ( .OUT(na1027_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1028_1),
                      .IN8(na2859_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1027_2 ( .OUT(na1027_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1027_1_i) );
// C_MX2b////      x92y81     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na433_1), .IN6(~na465_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x86y88     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1029_1 ( .OUT(na1029_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2860_1), .IN8(~na1030_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1029_2 ( .OUT(na1029_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1029_1_i) );
// C_MX2b////      x100y78     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na466_1), .IN6(~na434_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x85y88     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1031_1 ( .OUT(na1031_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2861_2), .IN8(~na1032_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1031_2 ( .OUT(na1031_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1031_1_i) );
// C_MX2b////      x94y76     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1032_1 ( .OUT(na1032_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na435_1), .IN6(~na467_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x85y91     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2862_1), .IN8(~na1034_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1033_2 ( .OUT(na1033_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1033_1_i) );
// C_MX2b////      x96y78     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1034_1 ( .OUT(na1034_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na436_2), .IN6(~na468_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x120y77     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_1 ( .OUT(na1035_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2691_1), .IN6(~na1036_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1035_2 ( .OUT(na1035_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1035_1_i) );
// C_MX2b////      x109y90     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1036_1 ( .OUT(na1036_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na437_2), .IN6(~na469_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x120y79     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1037_1 ( .OUT(na1037_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2697_1), .IN8(~na1038_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1037_2 ( .OUT(na1037_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1037_1_i) );
// C_MX2b////      x102y96     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1038_1 ( .OUT(na1038_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3017_2), .IN6(~na470_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x112y86     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2698_2), .IN8(~na1040_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1039_2 ( .OUT(na1039_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1039_1_i) );
// C_MX2b////      x114y84     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1040_1 ( .OUT(na1040_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na439_2), .IN8(~na471_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x116y79     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1041_1 ( .OUT(na1041_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2701_1), .IN8(~na1042_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1041_2 ( .OUT(na1041_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1041_1_i) );
// C_MX2b////      x108y78     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1042_1 ( .OUT(na1042_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na440_1), .IN6(~na3031_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x115y75     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1043_1 ( .OUT(na1043_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2702_2), .IN6(~na1044_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1043_2 ( .OUT(na1043_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1043_1_i) );
// C_MX2b////      x111y76     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1044_1 ( .OUT(na1044_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na473_2), .IN6(~na3018_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x111y85     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1045_1 ( .OUT(na1045_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2703_1), .IN6(~na1046_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1045_2 ( .OUT(na1045_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1045_1_i) );
// C_MX2b////      x111y78     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1046_1 ( .OUT(na1046_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na442_1), .IN8(~na474_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x116y78     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1047_1 ( .OUT(na1047_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2704_2), .IN8(~na1048_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1047_2 ( .OUT(na1047_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1047_1_i) );
// C_MX2b////      x108y74     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1048_1 ( .OUT(na1048_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na475_1), .IN6(~na443_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x121y76     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1049_1 ( .OUT(na1049_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2705_1), .IN6(~na1050_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1049_2 ( .OUT(na1049_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1049_1_i) );
// C_MX2b////      x111y72     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1050_1 ( .OUT(na1050_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na444_2), .IN6(~na476_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x122y88     80'h40_EC00_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_1 ( .OUT(na1051_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1052_1),
                      .IN8(na2731_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1051_2 ( .OUT(na1051_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1051_1_i) );
// C_MX2b////      x118y93     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1052_1 ( .OUT(na1052_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3035_2), .IN8(~na445_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x116y99     80'h40_EC00_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1053_1 ( .OUT(na1053_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1054_1),
                      .IN8(na2736_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1053_2 ( .OUT(na1053_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1053_1_i) );
// C_MX2b////      x118y97     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1054_1 ( .OUT(na1054_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na446_2), .IN6(~na3036_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x113y101     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_1 ( .OUT(na1055_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2737_2), .IN8(~na1056_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1055_2 ( .OUT(na1055_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1055_1_i) );
// C_MX2b////      x112y100     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1056_1 ( .OUT(na1056_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na447_1), .IN6(~na3037_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x111y94     80'h40_EC00_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1057_1 ( .OUT(na1057_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1058_1),
                      .IN8(na2740_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1057_2 ( .OUT(na1057_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1057_1_i) );
// C_MX2b////      x116y91     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1058_1 ( .OUT(na1058_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na448_2), .IN6(~na480_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x119y97     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_1 ( .OUT(na1059_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2741_2), .IN8(~na1060_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1059_2 ( .OUT(na1059_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1059_1_i) );
// C_MX2b////      x114y94     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1060_1 ( .OUT(na1060_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na481_2), .IN6(~na449_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x120y97     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_1 ( .OUT(na1061_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2742_1), .IN8(~na1062_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1061_2 ( .OUT(na1061_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1061_1_i) );
// C_MX2b////      x120y88     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1062_1 ( .OUT(na1062_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na450_1), .IN8(~na482_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x117y98     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_1 ( .OUT(na1063_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2743_2), .IN6(~na1064_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1063_2 ( .OUT(na1063_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1063_1_i) );
// C_MX2b////      x113y82     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na483_2), .IN6(~na451_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x116y100     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1065_1 ( .OUT(na1065_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2744_1), .IN8(~na1066_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1065_2 ( .OUT(na1065_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1065_1_i) );
// C_MX2b////      x118y98     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1066_1 ( .OUT(na1066_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3024_2), .IN6(~na484_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x115y104     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1067_1 ( .OUT(na1067_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2771_2), .IN8(~na1068_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1067_2 ( .OUT(na1067_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1067_1_i) );
// C_MX2b////      x108y96     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1068_1 ( .OUT(na1068_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na453_1), .IN8(~na3040_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x112y103     80'h40_EC00_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_1 ( .OUT(na1069_1_i), .IN1(1'b1), .IN2(~na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1070_1), .IN6(na2774_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1069_2 ( .OUT(na1069_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1069_1_i) );
// C_MX2b////      x105y99     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na454_2), .IN6(~na486_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x113y103     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_1 ( .OUT(na1071_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2775_1), .IN6(~na1072_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1071_2 ( .OUT(na1071_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1071_1_i) );
// C_MX2b////      x103y104     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1072_1 ( .OUT(na1072_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3025_2), .IN6(~na487_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x108y107     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1073_1 ( .OUT(na1073_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2778_2), .IN6(~na1074_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1073_2 ( .OUT(na1073_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1073_1_i) );
// C_MX2b////      x109y96     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1074_1 ( .OUT(na1074_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na456_2), .IN8(~na488_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x114y104     80'h40_EC00_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1075_1 ( .OUT(na1075_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2779_1), .IN6(~na1076_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1075_2 ( .OUT(na1075_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1075_1_i) );
// C_MX2b////      x107y98     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1076_1 ( .OUT(na1076_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na457_1), .IN6(~na3042_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x111y102     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1077_1 ( .OUT(na1077_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2780_2), .IN8(~na1078_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1077_2 ( .OUT(na1077_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1077_1_i) );
// C_MX2b////      x114y90     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1078_1 ( .OUT(na1078_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na490_1), .IN8(~na458_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x111y100     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_1 ( .OUT(na1079_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2781_1), .IN8(~na1080_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1079_2 ( .OUT(na1079_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1079_1_i) );
// C_MX2b////      x108y82     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1080_1 ( .OUT(na1080_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na491_2), .IN6(~na3028_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x112y104     80'h40_EC00_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1_i), .IN1(1'b1), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2782_2), .IN8(~na1082_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1081_2 ( .OUT(na1081_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1081_1_i) );
// C_MX2b////      x114y96     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1082_1 ( .OUT(na1082_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3029_2), .IN8(~na492_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x86y106     80'h40_EC00_00_0040_0C6A_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_1 ( .OUT(na1083_1_i), .IN1(1'b0), .IN2(~na1084_1), .IN3(1'b1), .IN4(na2904_2), .IN5(na1085_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na1083_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1083_2 ( .OUT(na1083_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1083_1_i) );
// C_MX4a/DST///      x83y108     80'h60_BC00_00_0040_0C9B_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1084_1 ( .OUT(na1084_1_i), .IN1(~na1085_1), .IN2(na3153_2), .IN3(1'b0), .IN4(~na2905_1), .IN5(1'b1), .IN6(na1084_1), .IN7(1'b1),
                      .IN8(~na1083_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0000)) 
           _a1084_2 ( .OUT(na1084_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1084_1_i) );
// C_AND/DST///      x87y105     80'h60_BC00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_1 ( .OUT(na1085_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1086_1), .IN8(na2906_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0000)) 
           _a1085_2 ( .OUT(na1085_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1085_1_i) );
// C_MX4b////      x84y109     80'h00_0018_00_0040_0A79_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1086_1 ( .OUT(na1086_1), .IN1(1'b1), .IN2(na3150_2), .IN3(na3152_2), .IN4(1'b1), .IN5(~na1085_1), .IN6(na2908_2), .IN7(na3215_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x99y87     80'h40_E418_00_0000_0888_F53F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_1 ( .OUT(na1087_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1010_1), .IN5(~na1087_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1087_5 ( .OUT(na1087_2), .CLK(1'b0), .EN(~na1103_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1087_1) );
// C_AND/D//AND/D      x98y91     80'h40_E400_80_0000_0C88_2F2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1089_1 ( .OUT(na1089_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1482_2), .IN8(~na1010_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1089_2 ( .OUT(na1089_1), .CLK(1'b0), .EN(~na1103_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1089_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1089_4 ( .OUT(na1089_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1482_1), .IN4(~na1010_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1089_5 ( .OUT(na1089_2), .CLK(1'b0), .EN(~na1103_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1089_2_i) );
// C_///AND/D      x99y92     80'h40_E400_80_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1090_4 ( .OUT(na1090_2_i), .IN1(~na3129_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1484_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1090_5 ( .OUT(na1090_2), .CLK(1'b0), .EN(~na1103_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1090_2_i) );
// C_MX4b////      x104y79     80'h00_0018_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1091_1 ( .OUT(na1091_1), .IN1(1'b1), .IN2(~na62_2), .IN3(1'b1), .IN4(~na1010_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1092_2),
                      .IN8(na1010_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y85     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1092_4 ( .OUT(na1092_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na66_1), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x103y93     80'h00_0018_00_0040_0C8B_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1094_1 ( .OUT(na1094_1), .IN1(na2909_1), .IN2(na3130_2), .IN3(1'b0), .IN4(~na429_1), .IN5(na1087_2), .IN6(1'b1), .IN7(~na2993_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x98y89     80'h00_0018_00_0000_0C88_DDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1095_1 ( .OUT(na1095_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3129_2), .IN6(na3160_2), .IN7(~na3155_2),
                      .IN8(na429_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y81     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1096_1 ( .OUT(na1096_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na2912_1), .IN7(na1103_2), .IN8(na3154_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x106y82     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1098_4 ( .OUT(na1098_2), .IN1(~na3129_2), .IN2(~na104_2), .IN3(1'b0), .IN4(~na1099_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y84     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1099_4 ( .OUT(na1099_2), .IN1(na1087_2), .IN2(na2855_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x102y95     80'h00_0018_00_0000_0C88_B3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1100_1 ( .OUT(na1100_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na3159_2), .IN7(na1103_2), .IN8(~na1010_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x101y96     80'h00_0018_00_0040_0C09_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1101_1 ( .OUT(na1101_1), .IN1(na1087_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1010_1), .IN5(1'b1), .IN6(~na62_2), .IN7(na1103_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y93     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1102_4 ( .OUT(na1102_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1103_1), .IN4(na1104_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x100y89     80'h00_0078_00_0000_0CEE_0B33
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1103_1 ( .OUT(na1103_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1087_1), .IN6(~na104_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1103_4 ( .OUT(na1103_2), .IN1(1'b0), .IN2(~na59_1), .IN3(1'b0), .IN4(~na1083_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x90y108     80'h00_0018_00_0040_0C0A_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1104_1 ( .OUT(na1104_1), .IN1(1'b0), .IN2(na1084_1), .IN3(1'b0), .IN4(na2918_2), .IN5(~na1085_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1083_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x102y84     80'h00_0018_00_0000_0888_EFAC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1105_1 ( .OUT(na1105_1), .IN1(1'b0), .IN2(na59_1), .IN3(na1103_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na1103_2), .IN8(na1010_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x98y95     80'h00_0018_00_0000_0888_EFEC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1106_1 ( .OUT(na1106_1), .IN1(1'b0), .IN2(na59_1), .IN3(na1103_2), .IN4(na3154_2), .IN5(1'b1), .IN6(1'b1), .IN7(na3151_2),
                      .IN8(na1010_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x93y100     80'h00_0060_00_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1107_4 ( .OUT(na1107_2), .IN1(na1087_2), .IN2(na2923_2), .IN3(1'b0), .IN4(~na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y92     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1108_1 ( .OUT(na1108_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1087_2), .IN6(na2855_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y96     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1109_1 ( .OUT(na1109_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2922_1), .IN7(na1103_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x96y87     80'h00_0018_00_0000_0888_5FE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1110_1 ( .OUT(na1110_1), .IN1(1'b0), .IN2(~na1108_1), .IN3(na66_1), .IN4(na429_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na66_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x107y81     80'h00_0018_00_0040_0C8A_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_1 ( .OUT(na1111_1), .IN1(1'b0), .IN2(na2923_1), .IN3(1'b0), .IN4(~na429_1), .IN5(~na1087_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na3217_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x106y83     80'h00_0018_00_0040_0C89_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1112_1 ( .OUT(na1112_1), .IN1(na3216_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na429_1), .IN5(na1087_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na3217_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x85y80     80'h00_0018_00_0040_0C05_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1113_1 ( .OUT(na1113_1), .IN1(na2925_1), .IN2(1'b0), .IN3(na2926_2), .IN4(1'b0), .IN5(1'b1), .IN6(na2348_2), .IN7(1'b1),
                      .IN8(na2350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x80y109     80'h00_EE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1114_1 ( .OUT(na1114_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2412_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2927_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1114_2 ( .OUT(na1114_1), .CLK(na1487_2), .EN(1'b1), .SR(na2404_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1114_1_i) );
// C_XOR////D      x97y87     80'hC0_EC18_00_0000_0666_AC0A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1115_1 ( .OUT(na1115_1), .IN1(na849_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na686_2), .IN7(na517_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1115_5 ( .OUT(na1115_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1115_1) );
// C_XOR/D///      x105y107     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_1 ( .OUT(na1116_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na518_1), .IN6(1'b0), .IN7(na685_1), .IN8(na899_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1116_2 ( .OUT(na1116_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1116_1_i) );
// C_///XOR/D      x104y106     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1117_4 ( .OUT(na1117_2_i), .IN1(1'b0), .IN2(na908_1), .IN3(na685_2), .IN4(na519_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1117_5 ( .OUT(na1117_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1117_2_i) );
// C_///XOR/D      x108y90     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1118_4 ( .OUT(na1118_2_i), .IN1(na688_1), .IN2(1'b0), .IN3(na912_1), .IN4(na520_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1118_5 ( .OUT(na1118_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1118_2_i) );
// C_XOR////D      x116y88     80'hC0_EC18_00_0000_0666_AAC5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1120_1 ( .OUT(na1120_1), .IN1(~na521_2), .IN2(1'b0), .IN3(1'b0), .IN4(na913_1), .IN5(na688_2), .IN6(1'b0), .IN7(na919_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1120_5 ( .OUT(na1120_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1120_1) );
// C_XOR////D      x117y68     80'hC0_EC18_00_0000_0666_C0AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_1 ( .OUT(na1121_1), .IN1(na921_1), .IN2(1'b0), .IN3(na690_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na522_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1121_5 ( .OUT(na1121_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1121_1) );
// C_///XOR/D      x110y68     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1122_4 ( .OUT(na1122_2_i), .IN1(na925_1), .IN2(1'b0), .IN3(na690_2), .IN4(na523_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1122_5 ( .OUT(na1122_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1122_2_i) );
// C_XOR/D///      x113y73     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1123_1 ( .OUT(na1123_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na927_1), .IN6(1'b0), .IN7(na3044_2), .IN8(na692_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1123_2 ( .OUT(na1123_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1123_1_i) );
// C_XOR////D      x81y110     80'hC0_EC18_00_0000_0666_0C0A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1124_1 ( .OUT(na1124_1), .IN1(na11_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na493_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1124_5 ( .OUT(na1124_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1124_1) );
// C_///XOR/D      x81y108     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1125_4 ( .OUT(na1125_2_i), .IN1(na430_2), .IN2(1'b0), .IN3(1'b0), .IN4(na69_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1125_5 ( .OUT(na1125_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1125_2_i) );
// C_XOR////D      x81y87     80'hC0_EC18_00_0000_0666_ACC5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1126_1 ( .OUT(na1126_1), .IN1(~na88_2), .IN2(1'b0), .IN3(1'b0), .IN4(na86_1), .IN5(1'b0), .IN6(na495_1), .IN7(na70_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1126_5 ( .OUT(na1126_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1126_1) );
// C_XOR////D      x85y74     80'hC0_EC18_00_0000_0666_0990
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1127_1 ( .OUT(na1127_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na95_1), .IN4(na86_1), .IN5(na88_2), .IN6(~na496_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1127_5 ( .OUT(na1127_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1127_1) );
// C_XOR////D      x86y65     80'hC0_EC18_00_0000_0666_A5C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1128_1 ( .OUT(na1128_1), .IN1(1'b0), .IN2(~na106_1), .IN3(1'b0), .IN4(na86_1), .IN5(~na497_2), .IN6(1'b0), .IN7(na95_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1128_5 ( .OUT(na1128_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1128_1) );
// C_XOR////D      x98y63     80'hC0_EC18_00_0000_0666_C50C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1), .IN1(1'b0), .IN2(na113_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na498_2), .IN6(1'b0), .IN7(1'b0), .IN8(na115_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1129_5 ( .OUT(na1129_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1129_1) );
// C_XOR////D      x85y64     80'hC0_EC18_00_0000_0666_C0CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1130_1 ( .OUT(na1130_1), .IN1(1'b0), .IN2(na113_1), .IN3(1'b0), .IN4(na499_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na122_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1130_5 ( .OUT(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1130_1) );
// C_XOR/D///      x88y66     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na500_1), .IN6(na2998_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1131_2 ( .OUT(na1131_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1131_1_i) );
// C_XOR////D      x112y99     80'hC0_EC18_00_0000_0666_A0A0
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1132_1 ( .OUT(na1132_1), .IN1(1'b0), .IN2(1'b0), .IN3(na693_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na501_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1132_5 ( .OUT(na1132_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1132_1) );
// C_///XOR/D      x107y103     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1133_4 ( .OUT(na1133_2_i), .IN1(na739_1), .IN2(1'b0), .IN3(na438_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1133_5 ( .OUT(na1133_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1133_2_i) );
// C_XOR////D      x117y78     80'hC0_EC18_00_0000_0666_3A3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1), .IN1(na749_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na752_2), .IN5(na750_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na503_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1134_5 ( .OUT(na1134_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1134_1) );
// C_XOR////D      x120y74     80'hC0_EC18_00_0000_0666_CA09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1), .IN1(na750_1), .IN2(~na755_1), .IN3(1'b0), .IN4(1'b0), .IN5(na504_2), .IN6(1'b0), .IN7(1'b0), .IN8(na752_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1135_5 ( .OUT(na1135_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1135_1) );
// C_XOR////D      x119y68     80'hC0_EC18_00_0000_0666_CC3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1136_1 ( .OUT(na1136_1), .IN1(na750_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na761_1), .IN5(1'b0), .IN6(na755_1), .IN7(1'b0), .IN8(na505_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1136_5 ( .OUT(na1136_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1136_1) );
// C_XOR/D///      x112y63     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na506_2), .IN7(na764_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1137_2 ( .OUT(na1137_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1137_1_i) );
// C_///XOR/D      x108y68     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1138_4 ( .OUT(na1138_2_i), .IN1(na769_1), .IN2(na507_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1138_5 ( .OUT(na1138_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1138_2_i) );
// C_XOR/D///      x112y68     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na771_1), .IN7(1'b0), .IN8(na508_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1139_2 ( .OUT(na1139_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1139_1_i) );
// C_XOR////D      x120y89     80'hC0_EC18_00_0000_0666_0A60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1), .IN1(1'b0), .IN2(1'b0), .IN3(na816_2), .IN4(na775_1), .IN5(na509_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1140_5 ( .OUT(na1140_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1140_1) );
// C_XOR////D      x117y80     80'hC0_EC18_00_0000_0666_0C0C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1), .IN1(1'b0), .IN2(na510_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na820_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1141_5 ( .OUT(na1141_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1141_1) );
// C_///XOR/D      x101y111     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1142_4 ( .OUT(na1142_2_i), .IN1(na829_1), .IN2(1'b0), .IN3(1'b0), .IN4(na511_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1142_5 ( .OUT(na1142_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1142_2_i) );
// C_XOR////D      x115y100     80'hC0_EC18_00_0000_0666_C05A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1143_1 ( .OUT(na1143_1), .IN1(na834_2), .IN2(1'b0), .IN3(~na512_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na775_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1143_5 ( .OUT(na1143_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1143_1) );
// C_XOR/D///      x106y110     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1144_1 ( .OUT(na1144_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na839_1), .IN6(1'b0), .IN7(na513_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1144_2 ( .OUT(na1144_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1144_1_i) );
// C_///XOR/D      x120y96     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1145_4 ( .OUT(na1145_2_i), .IN1(na842_1), .IN2(1'b0), .IN3(na450_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1145_5 ( .OUT(na1145_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1145_2_i) );
// C_XOR////D      x118y72     80'hC0_EC18_00_0000_0666_00AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1146_1 ( .OUT(na1146_1), .IN1(1'b0), .IN2(na515_2), .IN3(na845_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1146_5 ( .OUT(na1146_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1146_1) );
// C_XOR/D///      x109y108     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na847_1), .IN6(1'b0), .IN7(na452_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1147_2 ( .OUT(na1147_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1147_1_i) );
// C_///XOR/D      x89y111     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1148_4 ( .OUT(na1148_2_i), .IN1(1'b0), .IN2(na1124_1), .IN3(1'b0), .IN4(na525_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1148_5 ( .OUT(na1148_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1148_2_i) );
// C_XOR/D///      x81y108     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1149_1 ( .OUT(na1149_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na430_2), .IN6(1'b0), .IN7(na526_2), .IN8(na69_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1149_2 ( .OUT(na1149_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1149_1_i) );
// C_XOR/D///      x84y94     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1150_1 ( .OUT(na1150_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1126_1), .IN6(na527_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1150_2 ( .OUT(na1150_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1150_1_i) );
// C_///XOR/D      x88y75     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1151_4 ( .OUT(na1151_2_i), .IN1(1'b0), .IN2(na1127_1), .IN3(1'b0), .IN4(na528_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1151_5 ( .OUT(na1151_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1151_2_i) );
// C_XOR/D///      x90y65     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1152_1 ( .OUT(na1152_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1128_1), .IN8(na529_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1152_2 ( .OUT(na1152_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1152_1_i) );
// C_///XOR/D      x104y64     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1153_4 ( .OUT(na1153_2_i), .IN1(na530_1), .IN2(1'b0), .IN3(na1129_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1153_5 ( .OUT(na1153_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1153_2_i) );
// C_XOR/D///      x89y64     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_1 ( .OUT(na1154_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1130_1), .IN7(na531_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1154_2 ( .OUT(na1154_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1154_1_i) );
// C_XOR////D      x93y66     80'hC0_EC18_00_0000_0666_0ACA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_1 ( .OUT(na1155_1), .IN1(na128_1), .IN2(1'b0), .IN3(1'b0), .IN4(na532_2), .IN5(na500_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1155_5 ( .OUT(na1155_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1155_1) );
// C_///XOR/D      x111y98     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1156_4 ( .OUT(na1156_2_i), .IN1(1'b0), .IN2(na533_2), .IN3(na1132_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1156_5 ( .OUT(na1156_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1156_2_i) );
// C_///XOR/D      x110y107     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1157_4 ( .OUT(na1157_2_i), .IN1(na739_1), .IN2(1'b0), .IN3(na438_2), .IN4(na534_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1157_5 ( .OUT(na1157_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1157_2_i) );
// C_XOR/D///      x119y82     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1158_1 ( .OUT(na1158_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na535_1), .IN6(na1134_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1158_2 ( .OUT(na1158_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1158_1_i) );
// C_///XOR/D      x117y74     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1159_4 ( .OUT(na1159_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na536_2), .IN4(na1135_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1159_5 ( .OUT(na1159_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1159_2_i) );
// C_XOR/D///      x120y69     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1160_1 ( .OUT(na1160_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na537_1), .IN6(na1136_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1160_2 ( .OUT(na1160_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1160_1_i) );
// C_XOR////D      x111y64     80'hC0_EC18_00_0000_0666_0356
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_1 ( .OUT(na1161_1), .IN1(na765_1), .IN2(na766_1), .IN3(~na538_2), .IN4(1'b0), .IN5(1'b0), .IN6(~na506_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1161_5 ( .OUT(na1161_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1161_1) );
// C_XOR////D      x117y66     80'hC0_EC18_00_0000_0666_05A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1162_1 ( .OUT(na1162_1), .IN1(na765_1), .IN2(na507_1), .IN3(na744_1), .IN4(1'b0), .IN5(~na539_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1162_5 ( .OUT(na1162_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1162_1) );
// C_XOR////D      x120y66     80'hC0_EC18_00_0000_0666_0336
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_1 ( .OUT(na1163_1), .IN1(na765_1), .IN2(na772_2), .IN3(1'b0), .IN4(~na508_1), .IN5(1'b0), .IN6(~na540_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1163_5 ( .OUT(na1163_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1163_1) );
// C_///XOR/D      x119y89     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1164_4 ( .OUT(na1164_2_i), .IN1(na541_1), .IN2(1'b0), .IN3(na1140_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1164_5 ( .OUT(na1164_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1164_2_i) );
// C_XOR/D///      x115y78     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1141_1), .IN7(na542_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1165_2 ( .OUT(na1165_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1165_1_i) );
// C_XOR////D      x108y110     80'hC0_EC18_00_0000_0666_03C6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1166_1 ( .OUT(na1166_1), .IN1(na830_2), .IN2(na831_1), .IN3(1'b0), .IN4(na511_1), .IN5(1'b0), .IN6(~na543_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1166_5 ( .OUT(na1166_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1166_1) );
// C_///XOR/D      x123y102     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1167_4 ( .OUT(na1167_2_i), .IN1(1'b0), .IN2(na1143_1), .IN3(1'b0), .IN4(na544_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1167_5 ( .OUT(na1167_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1167_2_i) );
// C_XOR////D      x110y110     80'hC0_EC18_00_0000_0666_650A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1), .IN1(na834_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na545_1), .IN6(1'b0), .IN7(na513_2), .IN8(na840_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1168_5 ( .OUT(na1168_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1168_1) );
// C_///XOR/D      x120y94     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1169_4 ( .OUT(na1169_2_i), .IN1(na842_1), .IN2(1'b0), .IN3(na450_2), .IN4(na546_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1169_5 ( .OUT(na1169_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1169_2_i) );
// C_XOR/D///      x121y70     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_1 ( .OUT(na1170_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na547_1), .IN8(na1146_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1170_2 ( .OUT(na1170_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1170_1_i) );
// C_XOR/D///      x110y107     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_1 ( .OUT(na1171_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na847_1), .IN6(na548_2), .IN7(na452_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1171_2 ( .OUT(na1171_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1171_1_i) );
// C_///XOR/D      x100y88     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1172_4 ( .OUT(na1172_2_i), .IN1(na1115_1), .IN2(1'b0), .IN3(1'b0), .IN4(na549_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1172_5 ( .OUT(na1172_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1172_2_i) );
// C_XOR////D      x102y108     80'hC0_EC18_00_0000_0666_55CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_1 ( .OUT(na1173_1), .IN1(1'b0), .IN2(na550_2), .IN3(1'b0), .IN4(na899_1), .IN5(~na518_1), .IN6(1'b0), .IN7(~na685_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1173_5 ( .OUT(na1173_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1173_1) );
// C_XOR////D      x97y105     80'hC0_EC18_00_0000_0666_903C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1174_1 ( .OUT(na1174_1), .IN1(1'b0), .IN2(na908_1), .IN3(1'b0), .IN4(~na519_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na685_2), .IN8(na551_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1174_5 ( .OUT(na1174_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1174_1) );
// C_XOR////D      x113y96     80'hC0_EC18_00_0000_0666_6C3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1175_1 ( .OUT(na1175_1), .IN1(na688_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na520_2), .IN5(1'b0), .IN6(na552_1), .IN7(na850_1),
                      .IN8(na913_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1175_5 ( .OUT(na1175_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1175_1) );
// C_XOR/D///      x116y83     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1176_1 ( .OUT(na1176_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na553_1), .IN8(na1120_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1176_2 ( .OUT(na1176_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1176_1_i) );
// C_///XOR/D      x116y67     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1177_4 ( .OUT(na1177_2_i), .IN1(na554_2), .IN2(na1121_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1177_5 ( .OUT(na1177_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1177_2_i) );
// C_XOR////D      x110y65     80'hC0_EC18_00_0000_0666_3056
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1178_1 ( .OUT(na1178_1), .IN1(na925_1), .IN2(na555_2), .IN3(~na690_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(~na523_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1178_5 ( .OUT(na1178_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1178_1) );
// C_XOR////D      x104y73     80'hC0_EC18_00_0000_0666_3C3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1179_1 ( .OUT(na1179_1), .IN1(na927_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na692_2), .IN5(1'b0), .IN6(na556_2), .IN7(1'b0), .IN8(~na524_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1179_5 ( .OUT(na1179_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1179_1) );
// C_XOR/D///      x85y109     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1180_1 ( .OUT(na1180_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na557_1), .IN6(na1124_1), .IN7(1'b0), .IN8(na525_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1180_2 ( .OUT(na1180_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1180_1_i) );
// C_///XOR/D      x86y108     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1181_4 ( .OUT(na1181_2_i), .IN1(~na430_2), .IN2(na558_2), .IN3(~na526_2), .IN4(na69_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1181_5 ( .OUT(na1181_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1181_2_i) );
// C_XOR/D///      x87y94     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1182_1 ( .OUT(na1182_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1126_1), .IN6(na527_2), .IN7(na559_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1182_2 ( .OUT(na1182_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1182_1_i) );
// C_XOR/D///      x88y76     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1183_1 ( .OUT(na1183_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1127_1), .IN7(na560_1), .IN8(na528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1183_2 ( .OUT(na1183_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1183_1_i) );
// C_XOR/D///      x90y66     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1184_1 ( .OUT(na1184_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na561_1), .IN7(na1128_1), .IN8(na529_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1184_2 ( .OUT(na1184_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1184_1_i) );
// C_XOR/D///      x105y64     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1185_1 ( .OUT(na1185_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na530_1), .IN6(1'b0), .IN7(na1129_1), .IN8(na562_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1185_2 ( .OUT(na1185_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1185_1_i) );
// C_///XOR/D      x84y64     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1186_4 ( .OUT(na1186_2_i), .IN1(1'b0), .IN2(na1130_1), .IN3(na531_1), .IN4(na563_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1186_5 ( .OUT(na1186_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1186_2_i) );
// C_XOR/D///      x97y68     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1187_1 ( .OUT(na1187_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1155_1), .IN7(1'b0), .IN8(na564_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1187_2 ( .OUT(na1187_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1187_1_i) );
// C_///XOR/D      x111y104     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1188_4 ( .OUT(na1188_2_i), .IN1(1'b0), .IN2(na533_2), .IN3(na1132_1), .IN4(na565_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1188_5 ( .OUT(na1188_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1188_2_i) );
// C_XOR/D///      x105y101     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1189_1 ( .OUT(na1189_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na739_1), .IN6(na566_1), .IN7(~na438_2),
                      .IN8(~na534_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1189_2 ( .OUT(na1189_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1189_1_i) );
// C_///XOR/D      x120y83     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1190_4 ( .OUT(na1190_2_i), .IN1(na535_1), .IN2(na1134_1), .IN3(1'b0), .IN4(na567_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1190_5 ( .OUT(na1190_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1190_2_i) );
// C_XOR/D///      x117y74     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1191_1 ( .OUT(na1191_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na568_1), .IN7(na536_2), .IN8(na1135_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1191_2 ( .OUT(na1191_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1191_1_i) );
// C_XOR/D///      x119y70     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1192_1 ( .OUT(na1192_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na537_1), .IN6(na1136_1), .IN7(na569_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1192_2 ( .OUT(na1192_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1192_1_i) );
// C_///XOR/D      x112y63     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1193_4 ( .OUT(na1193_2_i), .IN1(na570_1), .IN2(na1161_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1193_5 ( .OUT(na1193_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1193_2_i) );
// C_XOR/D///      x115y68     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1194_1 ( .OUT(na1194_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1162_1), .IN7(1'b0), .IN8(na571_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1194_2 ( .OUT(na1194_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1194_1_i) );
// C_///XOR/D      x115y68     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1195_4 ( .OUT(na1195_2_i), .IN1(1'b0), .IN2(na572_2), .IN3(1'b0), .IN4(na1163_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1195_5 ( .OUT(na1195_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1195_2_i) );
// C_///XOR/D      x118y86     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1196_4 ( .OUT(na1196_2_i), .IN1(na541_1), .IN2(na573_1), .IN3(na1140_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1196_5 ( .OUT(na1196_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1196_2_i) );
// C_///XOR/D      x117y77     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1197_4 ( .OUT(na1197_2_i), .IN1(1'b0), .IN2(na1141_1), .IN3(na542_2), .IN4(na574_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1197_5 ( .OUT(na1197_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1197_2_i) );
// C_XOR/D///      x105y110     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1198_1 ( .OUT(na1198_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na575_1), .IN8(na1166_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1198_2 ( .OUT(na1198_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1198_1_i) );
// C_XOR/D///      x111y98     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_1 ( .OUT(na1199_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1143_1), .IN7(na576_2), .IN8(na544_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1199_2 ( .OUT(na1199_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1199_1_i) );
// C_///XOR/D      x107y108     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1200_4 ( .OUT(na1200_2_i), .IN1(1'b0), .IN2(na577_1), .IN3(1'b0), .IN4(na1168_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1200_5 ( .OUT(na1200_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1200_2_i) );
// C_///XOR/D      x118y94     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1201_4 ( .OUT(na1201_2_i), .IN1(na842_1), .IN2(na578_2), .IN3(~na450_2), .IN4(~na546_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1201_5 ( .OUT(na1201_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1201_2_i) );
// C_XOR/D///      x117y69     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1202_1 ( .OUT(na1202_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na579_1), .IN7(na547_1), .IN8(na1146_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1202_2 ( .OUT(na1202_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1202_1_i) );
// C_XOR/D///      x109y106     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1203_1 ( .OUT(na1203_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na847_1), .IN6(~na548_2), .IN7(~na452_2),
                      .IN8(na580_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1203_2 ( .OUT(na1203_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1203_1_i) );
// C_///XOR/D      x98y88     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1204_4 ( .OUT(na1204_2_i), .IN1(na1115_1), .IN2(na581_1), .IN3(1'b0), .IN4(na549_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1204_5 ( .OUT(na1204_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1204_2_i) );
// C_XOR/D///      x99y108     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1205_1 ( .OUT(na1205_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na582_2), .IN7(1'b0), .IN8(na1173_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1205_2 ( .OUT(na1205_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1205_1_i) );
// C_///XOR/D      x101y104     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1206_4 ( .OUT(na1206_2_i), .IN1(na1174_1), .IN2(na583_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1206_5 ( .OUT(na1206_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1206_2_i) );
// C_XOR/D///      x117y93     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1207_1 ( .OUT(na1207_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1175_1), .IN7(1'b0), .IN8(na584_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1207_2 ( .OUT(na1207_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1207_1_i) );
// C_///XOR/D      x119y85     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1208_4 ( .OUT(na1208_2_i), .IN1(1'b0), .IN2(na585_1), .IN3(na553_1), .IN4(na1120_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1208_5 ( .OUT(na1208_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1208_2_i) );
// C_///XOR/D      x114y64     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1209_4 ( .OUT(na1209_2_i), .IN1(na554_2), .IN2(na1121_1), .IN3(na586_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1209_5 ( .OUT(na1209_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1209_2_i) );
// C_///XOR/D      x101y66     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1210_4 ( .OUT(na1210_2_i), .IN1(1'b0), .IN2(na587_1), .IN3(na1178_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1210_5 ( .OUT(na1210_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1210_2_i) );
// C_XOR/D///      x110y68     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1211_1 ( .OUT(na1211_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1179_1), .IN8(na588_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1211_2 ( .OUT(na1211_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1211_1_i) );
// C_///XOR/D      x88y106     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1212_4 ( .OUT(na1212_2_i), .IN1(~na557_1), .IN2(na1124_1), .IN3(na428_1), .IN4(~na525_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1212_5 ( .OUT(na1212_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1212_2_i) );
// C_XOR/D///      x82y108     80'hC0_EC00_00_0000_0666_59CA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1213_1 ( .OUT(na1213_1_i), .IN1(na430_1), .IN2(1'b0), .IN3(1'b0), .IN4(na69_1), .IN5(~na430_2), .IN6(na558_2), .IN7(~na526_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1213_2 ( .OUT(na1213_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1213_1_i) );
// C_XOR/D///      x88y91     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1214_1 ( .OUT(na1214_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1126_1), .IN6(na431_1), .IN7(~na559_1),
                      .IN8(~na3045_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1214_2 ( .OUT(na1214_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1214_1_i) );
// C_XOR/D///      x89y78     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1215_1 ( .OUT(na1215_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na432_2), .IN6(na1127_1), .IN7(~na560_1),
                      .IN8(~na528_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1215_2 ( .OUT(na1215_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1215_1_i) );
// C_XOR/D///      x92y69     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1216_1 ( .OUT(na1216_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na433_1), .IN6(~na561_1), .IN7(na1128_1),
                      .IN8(~na529_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1216_2 ( .OUT(na1216_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1216_1_i) );
// C_///XOR/D      x101y65     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1217_4 ( .OUT(na1217_2_i), .IN1(~na530_1), .IN2(na434_2), .IN3(na1129_1), .IN4(~na562_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1217_5 ( .OUT(na1217_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1217_2_i) );
// C_XOR/D///      x95y65     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1218_1 ( .OUT(na1218_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na435_1), .IN6(na1130_1), .IN7(~na531_1),
                      .IN8(~na563_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1218_2 ( .OUT(na1218_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1218_1_i) );
// C_XOR/D///      x99y65     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1219_1 ( .OUT(na1219_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na436_2), .IN6(na1155_1), .IN7(1'b0), .IN8(na564_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1219_2 ( .OUT(na1219_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1219_1_i) );
// C_///XOR/D      x105y101     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1220_4 ( .OUT(na1220_2_i), .IN1(na437_2), .IN2(~na533_2), .IN3(na1132_1), .IN4(~na565_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1220_5 ( .OUT(na1220_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1220_2_i) );
// C_XOR/D///      x106y102     80'hC0_EC00_00_0000_0666_60A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1221_1 ( .OUT(na1221_1_i), .IN1(na739_1), .IN2(na566_1), .IN3(na438_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na438_2),
                      .IN8(~na534_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1221_2 ( .OUT(na1221_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1221_1_i) );
// C_XOR/D///      x118y82     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1222_1 ( .OUT(na1222_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na535_1), .IN6(na1134_1), .IN7(na439_2),
                      .IN8(~na567_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1222_2 ( .OUT(na1222_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1222_1_i) );
// C_///XOR/D      x119y82     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1223_4 ( .OUT(na1223_2_i), .IN1(na440_1), .IN2(~na568_1), .IN3(~na536_2), .IN4(na1135_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1223_5 ( .OUT(na1223_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1223_2_i) );
// C_///XOR/D      x117y71     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1224_4 ( .OUT(na1224_2_i), .IN1(~na537_1), .IN2(na1136_1), .IN3(~na569_1), .IN4(na441_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1224_5 ( .OUT(na1224_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1224_2_i) );
// C_///XOR/D      x111y67     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1225_4 ( .OUT(na1225_2_i), .IN1(na570_1), .IN2(na1161_1), .IN3(na442_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1225_5 ( .OUT(na1225_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1225_2_i) );
// C_XOR/D///      x111y70     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1226_1 ( .OUT(na1226_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3019_2), .IN6(na1162_1), .IN7(1'b0), .IN8(na571_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1226_2 ( .OUT(na1226_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1226_1_i) );
// C_XOR/D///      x113y71     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1227_1 ( .OUT(na1227_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na444_2), .IN6(na572_2), .IN7(1'b0), .IN8(na1163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1227_2 ( .OUT(na1227_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1227_1_i) );
// C_///XOR/D      x120y87     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1228_4 ( .OUT(na1228_2_i), .IN1(~na541_1), .IN2(~na573_1), .IN3(na1140_1), .IN4(na445_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1228_5 ( .OUT(na1228_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1228_2_i) );
// C_XOR/D///      x114y80     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1229_1 ( .OUT(na1229_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na446_2), .IN6(na1141_1), .IN7(~na542_2),
                      .IN8(~na574_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1229_2 ( .OUT(na1229_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1229_1_i) );
// C_XOR/D///      x105y108     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1230_1 ( .OUT(na1230_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na447_1), .IN6(1'b0), .IN7(na575_1), .IN8(na1166_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1230_2 ( .OUT(na1230_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1230_1_i) );
// C_///XOR/D      x115y98     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1231_4 ( .OUT(na1231_2_i), .IN1(na448_2), .IN2(na1143_1), .IN3(~na576_2), .IN4(~na544_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1231_5 ( .OUT(na1231_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1231_2_i) );
// C_///XOR/D      x109y108     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1232_4 ( .OUT(na1232_2_i), .IN1(na3050_2), .IN2(na449_1), .IN3(1'b0), .IN4(na1168_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1232_5 ( .OUT(na1232_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1232_2_i) );
// C_XOR/D///      x120y92     80'hC0_EC00_00_0000_0666_5C9A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1233_1 ( .OUT(na1233_1_i), .IN1(na842_1), .IN2(1'b0), .IN3(na450_1), .IN4(~na546_1), .IN5(1'b0), .IN6(na578_2), .IN7(~na450_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1233_2 ( .OUT(na1233_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1233_1_i) );
// C_XOR/D///      x117y72     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1234_1 ( .OUT(na1234_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3051_2), .IN6(na451_1), .IN7(~na547_1),
                      .IN8(na1146_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1234_2 ( .OUT(na1234_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1234_1_i) );
// C_XOR/D///      x110y106     80'hC0_EC00_00_0000_0666_5069
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1235_1 ( .OUT(na1235_1_i), .IN1(na847_1), .IN2(~na548_2), .IN3(na452_1), .IN4(na580_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na452_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1235_2 ( .OUT(na1235_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1235_1_i) );
// C_///XOR/D      x98y90     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1236_4 ( .OUT(na1236_2_i), .IN1(na1115_1), .IN2(~na581_1), .IN3(na453_1), .IN4(~na549_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1236_5 ( .OUT(na1236_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1236_2_i) );
// C_XOR/D///      x102y107     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1237_1 ( .OUT(na1237_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na454_2), .IN6(na582_2), .IN7(1'b0), .IN8(na1173_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1237_2 ( .OUT(na1237_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1237_1_i) );
// C_XOR/D///      x101y106     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1238_1 ( .OUT(na1238_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1174_1), .IN6(na583_1), .IN7(na455_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1238_2 ( .OUT(na1238_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1238_1_i) );
// C_XOR/D///      x109y92     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_1 ( .OUT(na1239_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1175_1), .IN7(na456_2), .IN8(na584_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1239_2 ( .OUT(na1239_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1239_1_i) );
// C_XOR/D///      x117y86     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1240_1 ( .OUT(na1240_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na457_1), .IN6(~na585_1), .IN7(~na553_1),
                      .IN8(na1120_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1240_2 ( .OUT(na1240_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1240_1_i) );
// C_XOR/D///      x110y72     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1241_1 ( .OUT(na1241_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na554_2), .IN6(na1121_1), .IN7(~na586_2),
                      .IN8(na458_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1241_2 ( .OUT(na1241_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1241_1_i) );
// C_///XOR/D      x107y68     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1242_4 ( .OUT(na1242_2_i), .IN1(na459_2), .IN2(na587_1), .IN3(na1178_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1242_5 ( .OUT(na1242_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1242_2_i) );
// C_XOR/D///      x112y73     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1243_1 ( .OUT(na1243_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na460_2), .IN6(1'b0), .IN7(na1179_1), .IN8(na588_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1243_2 ( .OUT(na1243_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1243_1_i) );
// C_XOR////D      x83y109     80'hC0_EC18_00_0000_0666_0A0A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1244_1 ( .OUT(na1244_1), .IN1(na11_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na589_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1244_5 ( .OUT(na1244_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1244_1) );
// C_///XOR/D      x83y105     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1245_4 ( .OUT(na1245_2_i), .IN1(1'b0), .IN2(na470_2), .IN3(1'b0), .IN4(na69_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1245_5 ( .OUT(na1245_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1245_2_i) );
// C_XOR////D      x82y87     80'hC0_EC18_00_0000_0666_C560
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1246_1 ( .OUT(na1246_1), .IN1(1'b0), .IN2(1'b0), .IN3(na70_1), .IN4(na86_1), .IN5(~na88_2), .IN6(1'b0), .IN7(1'b0), .IN8(na591_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1246_5 ( .OUT(na1246_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1246_1) );
// C_XOR////D      x85y76     80'hC0_EC18_00_0000_0666_059A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1247_1 ( .OUT(na1247_1), .IN1(na88_2), .IN2(1'b0), .IN3(~na95_1), .IN4(na86_1), .IN5(~na592_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1247_5 ( .OUT(na1247_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1247_1) );
// C_XOR////D      x87y66     80'hC0_EC18_00_0000_0666_0363
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1248_1 ( .OUT(na1248_1), .IN1(1'b0), .IN2(~na106_1), .IN3(na95_1), .IN4(na86_1), .IN5(1'b0), .IN6(~na593_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1248_5 ( .OUT(na1248_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1248_1) );
// C_XOR////D      x95y64     80'hC0_EC18_00_0000_0666_03CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1249_1 ( .OUT(na1249_1), .IN1(1'b0), .IN2(na113_1), .IN3(1'b0), .IN4(na115_1), .IN5(1'b0), .IN6(~na594_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1249_5 ( .OUT(na1249_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1249_1) );
// C_XOR////D      x87y64     80'hC0_EC18_00_0000_0666_006C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1250_1 ( .OUT(na1250_1), .IN1(1'b0), .IN2(na113_1), .IN3(na595_2), .IN4(na122_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1250_5 ( .OUT(na1250_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1250_1) );
// C_XOR/D///      x90y67     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1251_1 ( .OUT(na1251_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na128_1), .IN6(1'b0), .IN7(na596_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1251_2 ( .OUT(na1251_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1251_1_i) );
// C_XOR////D      x120y95     80'hC0_EC18_00_0000_0666_00AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1252_1 ( .OUT(na1252_1), .IN1(na597_2), .IN2(1'b0), .IN3(na693_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1252_5 ( .OUT(na1252_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1252_1) );
// C_///XOR/D      x108y103     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1253_4 ( .OUT(na1253_2_i), .IN1(na739_1), .IN2(1'b0), .IN3(1'b0), .IN4(na478_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1253_5 ( .OUT(na1253_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1253_2_i) );
// C_XOR////D      x119y78     80'hC0_EC18_00_0000_0666_0A6A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1254_1 ( .OUT(na1254_1), .IN1(na750_1), .IN2(1'b0), .IN3(~na599_1), .IN4(~na752_2), .IN5(na749_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1254_5 ( .OUT(na1254_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1254_1) );
// C_XOR////D      x120y71     80'hC0_EC18_00_0000_0666_C0A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1255_1 ( .OUT(na1255_1), .IN1(na750_1), .IN2(~na755_1), .IN3(na600_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na752_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1255_5 ( .OUT(na1255_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1255_1) );
// C_XOR////D      x120y68     80'hC0_EC18_00_0000_0666_0096
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1256_1 ( .OUT(na1256_1), .IN1(na750_1), .IN2(na755_1), .IN3(na601_1), .IN4(~na761_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1256_5 ( .OUT(na1256_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1256_1) );
// C_XOR/D///      x114y64     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1257_1 ( .OUT(na1257_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na602_2), .IN6(1'b0), .IN7(na764_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1257_2 ( .OUT(na1257_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1257_1_i) );
// C_///XOR/D      x109y66     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1258_4 ( .OUT(na1258_2_i), .IN1(na769_1), .IN2(1'b0), .IN3(1'b0), .IN4(na603_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1258_5 ( .OUT(na1258_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1258_2_i) );
// C_XOR/D///      x113y67     80'hC0_EC00_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1259_1 ( .OUT(na1259_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na771_1), .IN7(na604_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1259_2 ( .OUT(na1259_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1259_1_i) );
// C_XOR////D      x116y87     80'hC0_EC18_00_0000_0666_0C60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1260_1 ( .OUT(na1260_1), .IN1(1'b0), .IN2(1'b0), .IN3(na816_2), .IN4(na775_1), .IN5(1'b0), .IN6(na605_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1260_5 ( .OUT(na1260_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1260_1) );
// C_XOR////D      x116y75     80'hC0_EC18_00_0000_0666_00CC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1261_1 ( .OUT(na1261_1), .IN1(1'b0), .IN2(na820_1), .IN3(1'b0), .IN4(na606_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1261_5 ( .OUT(na1261_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1261_1) );
// C_///XOR/D      x100y111     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1262_4 ( .OUT(na1262_2_i), .IN1(na829_1), .IN2(na607_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1262_5 ( .OUT(na1262_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1262_2_i) );
// C_XOR////D      x114y99     80'hC0_EC18_00_0000_0666_05CA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1263_1 ( .OUT(na1263_1), .IN1(na834_2), .IN2(1'b0), .IN3(1'b0), .IN4(na775_1), .IN5(~na608_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1263_5 ( .OUT(na1263_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1263_1) );
// C_XOR/D///      x103y110     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1264_1 ( .OUT(na1264_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na839_1), .IN6(na609_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1264_2 ( .OUT(na1264_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1264_1_i) );
// C_///XOR/D      x119y98     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1265_4 ( .OUT(na1265_2_i), .IN1(na842_1), .IN2(1'b0), .IN3(na490_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1265_5 ( .OUT(na1265_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1265_2_i) );
// C_XOR////D      x119y74     80'hC0_EC18_00_0000_0666_0060
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1266_1 ( .OUT(na1266_1), .IN1(1'b0), .IN2(1'b0), .IN3(na845_1), .IN4(na611_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1266_5 ( .OUT(na1266_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1266_1) );
// C_XOR/D///      x113y104     80'hC0_EC00_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1267_1 ( .OUT(na1267_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na847_1), .IN6(1'b0), .IN7(1'b0), .IN8(na492_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1267_2 ( .OUT(na1267_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1267_1_i) );
// C_///XOR/D      x90y105     80'hC0_EC00_80_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1268_4 ( .OUT(na1268_2_i), .IN1(na849_1), .IN2(1'b0), .IN3(1'b0), .IN4(na461_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1268_5 ( .OUT(na1268_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1268_2_i) );
// C_XOR/D///      x97y110     80'hC0_EC00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1269_1 ( .OUT(na1269_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na462_2), .IN7(1'b0), .IN8(na899_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1269_2 ( .OUT(na1269_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1269_1_i) );
// C_XOR////D      x89y109     80'hC0_EC18_00_0000_0666_00AC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1270_1 ( .OUT(na1270_1), .IN1(1'b0), .IN2(na908_1), .IN3(na615_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1270_5 ( .OUT(na1270_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1270_1) );
// C_XOR////D      x108y101     80'hC0_EC18_00_0000_0666_0360
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_1 ( .OUT(na1271_1), .IN1(1'b0), .IN2(1'b0), .IN3(na850_1), .IN4(na913_1), .IN5(1'b0), .IN6(~na616_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1271_5 ( .OUT(na1271_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1271_1) );
// C_///XOR/D      x106y89     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1272_4 ( .OUT(na1272_2_i), .IN1(1'b0), .IN2(na617_1), .IN3(na918_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1272_5 ( .OUT(na1272_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1272_2_i) );
// C_XOR////D      x115y67     80'hC0_EC18_00_0000_0666_00AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1273_1 ( .OUT(na1273_1), .IN1(na921_1), .IN2(1'b0), .IN3(na618_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1273_5 ( .OUT(na1273_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1273_1) );
// C_XOR/D///      x104y68     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1274_1 ( .OUT(na1274_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na925_1), .IN6(na467_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1274_2 ( .OUT(na1274_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1274_1_i) );
// C_///XOR/D      x106y78     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1275_4 ( .OUT(na1275_2_i), .IN1(na927_1), .IN2(na468_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1275_5 ( .OUT(na1275_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1275_2_i) );
// C_XOR/D///      x86y110     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1276_1 ( .OUT(na1276_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1244_1), .IN6(1'b0), .IN7(na621_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1276_2 ( .OUT(na1276_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1276_1_i) );
// C_///XOR/D      x84y107     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1277_4 ( .OUT(na1277_2_i), .IN1(1'b0), .IN2(na470_2), .IN3(na622_2), .IN4(na69_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1277_5 ( .OUT(na1277_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1277_2_i) );
// C_///XOR/D      x84y94     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1278_4 ( .OUT(na1278_2_i), .IN1(na623_1), .IN2(1'b0), .IN3(na1246_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1278_5 ( .OUT(na1278_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1278_2_i) );
// C_XOR/D///      x86y76     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1279_1 ( .OUT(na1279_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na624_2), .IN6(na1247_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1279_2 ( .OUT(na1279_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1279_1_i) );
// C_///XOR/D      x83y67     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1280_4 ( .OUT(na1280_2_i), .IN1(1'b0), .IN2(na1248_1), .IN3(1'b0), .IN4(na625_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1280_5 ( .OUT(na1280_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1280_2_i) );
// C_XOR/D///      x104y64     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1281_1 ( .OUT(na1281_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na626_2), .IN6(na1249_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1281_2 ( .OUT(na1281_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1281_1_i) );
// C_///XOR/D      x95y65     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1282_4 ( .OUT(na1282_2_i), .IN1(1'b0), .IN2(na1250_1), .IN3(1'b0), .IN4(na627_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1282_5 ( .OUT(na1282_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1282_2_i) );
// C_XOR////D      x92y65     80'hC0_EC18_00_0000_0666_00A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1283_1 ( .OUT(na1283_1), .IN1(na128_1), .IN2(na628_1), .IN3(na596_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1283_5 ( .OUT(na1283_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1283_1) );
// C_XOR/D///      x121y96     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1284_1 ( .OUT(na1284_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na629_2), .IN6(1'b0), .IN7(na1252_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1284_2 ( .OUT(na1284_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1284_1_i) );
// C_///XOR/D      x109y106     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1285_4 ( .OUT(na1285_2_i), .IN1(na739_1), .IN2(1'b0), .IN3(na630_1), .IN4(na478_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1285_5 ( .OUT(na1285_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1285_2_i) );
// C_///XOR/D      x123y84     80'hC0_EC00_80_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1286_4 ( .OUT(na1286_2_i), .IN1(na631_1), .IN2(na1254_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1286_5 ( .OUT(na1286_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1286_2_i) );
// C_XOR/D///      x121y74     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1287_1 ( .OUT(na1287_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1255_1), .IN8(na632_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1287_2 ( .OUT(na1287_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1287_1_i) );
// C_///XOR/D      x121y69     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1288_4 ( .OUT(na1288_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na633_2), .IN4(na1256_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1288_5 ( .OUT(na1288_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1288_2_i) );
// C_XOR////D      x112y65     80'hC0_EC18_00_0000_0666_0536
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_1 ( .OUT(na1289_1), .IN1(na765_1), .IN2(na766_1), .IN3(1'b0), .IN4(~na634_1), .IN5(~na602_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1289_5 ( .OUT(na1289_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1289_1) );
// C_XOR////D      x118y66     80'hC0_EC18_00_0000_0666_036A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1290_1 ( .OUT(na1290_1), .IN1(na765_1), .IN2(1'b0), .IN3(na744_1), .IN4(na603_1), .IN5(1'b0), .IN6(~na635_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1290_5 ( .OUT(na1290_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1290_1) );
// C_XOR////D      x120y67     80'hC0_EC18_00_0000_0666_0066
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1291_1 ( .OUT(na1291_1), .IN1(na765_1), .IN2(na772_2), .IN3(~na604_2), .IN4(~na636_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1291_5 ( .OUT(na1291_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1291_1) );
// C_XOR/D///      x120y83     80'hC0_EC00_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1292_1 ( .OUT(na1292_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1260_1), .IN8(na637_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1292_2 ( .OUT(na1292_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1292_1_i) );
// C_///XOR/D      x116y74     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1293_4 ( .OUT(na1293_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1261_1), .IN4(na638_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1293_5 ( .OUT(na1293_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1293_2_i) );
// C_XOR////D      x104y110     80'hC0_EC18_00_0000_0666_0906
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1294_1 ( .OUT(na1294_1), .IN1(na830_2), .IN2(na831_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na639_2), .IN6(na607_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1294_5 ( .OUT(na1294_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1294_1) );
// C_XOR/D///      x115y98     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1295_1 ( .OUT(na1295_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na640_1), .IN6(1'b0), .IN7(na1263_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1295_2 ( .OUT(na1295_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1295_1_i) );
// C_XOR////D      x109y110     80'hC0_EC18_00_0000_0666_C056
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1296_1 ( .OUT(na1296_1), .IN1(na834_2), .IN2(na609_1), .IN3(~na641_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na840_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1296_5 ( .OUT(na1296_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1296_1) );
// C_XOR/D///      x120y94     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1297_1 ( .OUT(na1297_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na842_1), .IN6(1'b0), .IN7(na490_2), .IN8(na642_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1297_2 ( .OUT(na1297_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1297_1_i) );
// C_///XOR/D      x120y69     80'hC0_EC00_80_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1298_4 ( .OUT(na1298_2_i), .IN1(1'b0), .IN2(na1266_1), .IN3(1'b0), .IN4(na643_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1298_5 ( .OUT(na1298_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1298_2_i) );
// C_///XOR/D      x112y107     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1299_4 ( .OUT(na1299_2_i), .IN1(na847_1), .IN2(1'b0), .IN3(na644_1), .IN4(na492_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1299_5 ( .OUT(na1299_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1299_2_i) );
// C_XOR/D///      x87y99     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1300_1 ( .OUT(na1300_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na849_1), .IN6(1'b0), .IN7(na645_2), .IN8(na461_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1300_2 ( .OUT(na1300_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1300_1_i) );
// C_///XOR/D      x96y109     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1301_4 ( .OUT(na1301_2_i), .IN1(na646_1), .IN2(na462_2), .IN3(1'b0), .IN4(na899_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1301_5 ( .OUT(na1301_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1301_2_i) );
// C_XOR/D///      x89y108     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1302_1 ( .OUT(na1302_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1270_1), .IN6(1'b0), .IN7(na647_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1302_2 ( .OUT(na1302_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1302_1_i) );
// C_///XOR/D      x106y103     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1303_4 ( .OUT(na1303_2_i), .IN1(na648_1), .IN2(1'b0), .IN3(na1271_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1303_5 ( .OUT(na1303_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1303_2_i) );
// C_XOR////D      x115y91     80'hC0_EC18_00_0000_0666_306C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1304_1 ( .OUT(na1304_1), .IN1(1'b0), .IN2(na617_1), .IN3(na919_2), .IN4(na913_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(~na649_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1304_5 ( .OUT(na1304_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1304_1) );
// C_XOR/D///      x113y66     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1305_1 ( .OUT(na1305_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1273_1), .IN6(na650_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1305_2 ( .OUT(na1305_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1305_1_i) );
// C_XOR/D///      x106y67     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1306_1 ( .OUT(na1306_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na651_2), .IN6(na467_2), .IN7(1'b0), .IN8(na3128_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1306_2 ( .OUT(na1306_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1306_1_i) );
// C_///XOR/D      x107y78     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1307_4 ( .OUT(na1307_2_i), .IN1(na927_1), .IN2(na468_2), .IN3(1'b0), .IN4(na652_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1307_5 ( .OUT(na1307_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1307_2_i) );
// C_XOR/D///      x87y112     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_1 ( .OUT(na1308_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1244_1), .IN6(1'b0), .IN7(na621_1), .IN8(na653_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1308_2 ( .OUT(na1308_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1308_1_i) );
// C_XOR/D///      x83y106     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1309_1 ( .OUT(na1309_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na654_1), .IN6(~na470_2), .IN7(~na622_2),
                      .IN8(na69_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1309_2 ( .OUT(na1309_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1309_1_i) );
// C_XOR/D///      x86y91     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1310_1 ( .OUT(na1310_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na623_1), .IN6(na655_2), .IN7(na1246_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1310_2 ( .OUT(na1310_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1310_1_i) );
// C_///XOR/D      x89y78     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1311_4 ( .OUT(na1311_2_i), .IN1(na624_2), .IN2(na1247_1), .IN3(na656_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1311_5 ( .OUT(na1311_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1311_2_i) );
// C_///XOR/D      x88y66     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1312_4 ( .OUT(na1312_2_i), .IN1(1'b0), .IN2(na1248_1), .IN3(na657_2), .IN4(na625_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1312_5 ( .OUT(na1312_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1312_2_i) );
// C_XOR/D///      x100y64     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na626_2), .IN6(na1249_1), .IN7(1'b0), .IN8(na658_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1313_2 ( .OUT(na1313_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1313_1_i) );
// C_XOR/D///      x92y64     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1314_1 ( .OUT(na1314_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1250_1), .IN7(na659_2), .IN8(na627_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1314_2 ( .OUT(na1314_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1314_1_i) );
// C_///XOR/D      x93y68     80'hC0_EC00_80_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1315_4 ( .OUT(na1315_2_i), .IN1(1'b0), .IN2(na660_1), .IN3(na1283_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1315_5 ( .OUT(na1315_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1315_2_i) );
// C_XOR/D///      x119y96     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1316_1 ( .OUT(na1316_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na629_2), .IN6(1'b0), .IN7(na1252_1), .IN8(na661_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1316_2 ( .OUT(na1316_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1316_1_i) );
// C_///XOR/D      x112y106     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1317_4 ( .OUT(na1317_2_i), .IN1(na739_1), .IN2(na662_1), .IN3(~na630_1), .IN4(~na478_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1317_5 ( .OUT(na1317_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1317_2_i) );
// C_XOR/D///      x120y85     80'hC0_EC00_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1318_1 ( .OUT(na1318_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na631_1), .IN6(na1254_1), .IN7(1'b0), .IN8(na663_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1318_2 ( .OUT(na1318_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1318_1_i) );
// C_///XOR/D      x119y71     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1319_4 ( .OUT(na1319_2_i), .IN1(1'b0), .IN2(na664_1), .IN3(na1255_1), .IN4(na632_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1319_5 ( .OUT(na1319_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1319_2_i) );
// C_///XOR/D      x119y72     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1320_4 ( .OUT(na1320_2_i), .IN1(1'b0), .IN2(na665_2), .IN3(na633_2), .IN4(na1256_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1320_5 ( .OUT(na1320_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1320_2_i) );
// C_XOR/D///      x120y65     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1321_1 ( .OUT(na1321_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na666_1), .IN6(1'b0), .IN7(na1289_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1321_2 ( .OUT(na1321_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1321_1_i) );
// C_///XOR/D      x113y68     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1322_4 ( .OUT(na1322_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na667_2), .IN4(na1290_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1322_5 ( .OUT(na1322_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1322_2_i) );
// C_XOR/D///      x116y69     80'hC0_EC00_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_1 ( .OUT(na1323_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na668_1), .IN6(1'b0), .IN7(na1291_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1323_2 ( .OUT(na1323_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1323_1_i) );
// C_///XOR/D      x120y85     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1324_4 ( .OUT(na1324_2_i), .IN1(na669_2), .IN2(1'b0), .IN3(na1260_1), .IN4(na637_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1324_5 ( .OUT(na1324_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1324_2_i) );
// C_///XOR/D      x116y77     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1325_4 ( .OUT(na1325_2_i), .IN1(1'b0), .IN2(na670_1), .IN3(na1261_1), .IN4(na638_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1325_5 ( .OUT(na1325_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1325_2_i) );
// C_///XOR/D      x103y110     80'hC0_EC00_80_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1326_4 ( .OUT(na1326_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(na671_2), .IN4(na1294_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1326_5 ( .OUT(na1326_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1326_2_i) );
// C_///XOR/D      x120y98     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1327_4 ( .OUT(na1327_2_i), .IN1(na640_1), .IN2(na672_1), .IN3(na1263_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1327_5 ( .OUT(na1327_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1327_2_i) );
// C_XOR/D///      x107y109     80'hC0_EC00_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1328_1 ( .OUT(na1328_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na673_2), .IN6(na1296_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1328_2 ( .OUT(na1328_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1328_1_i) );
// C_XOR/D///      x122y93     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1329_1 ( .OUT(na1329_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na842_1), .IN6(na674_1), .IN7(~na490_2),
                      .IN8(~na642_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1329_2 ( .OUT(na1329_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1329_1_i) );
// C_XOR/D///      x119y71     80'hC0_EC00_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1330_1 ( .OUT(na1330_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1266_1), .IN7(na675_2), .IN8(na643_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1330_2 ( .OUT(na1330_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1330_1_i) );
// C_///XOR/D      x111y103     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1331_4 ( .OUT(na1331_2_i), .IN1(na847_1), .IN2(na676_1), .IN3(~na644_1), .IN4(~na492_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1331_5 ( .OUT(na1331_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1331_2_i) );
// C_///XOR/D      x90y103     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1332_4 ( .OUT(na1332_2_i), .IN1(na849_1), .IN2(na677_2), .IN3(~na645_2), .IN4(~na461_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1332_5 ( .OUT(na1332_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1332_2_i) );
// C_XOR/D///      x97y109     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na646_1), .IN6(~na462_2), .IN7(na678_1),
                      .IN8(na899_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1333_2 ( .OUT(na1333_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1333_1_i) );
// C_XOR/D///      x90y105     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1334_1 ( .OUT(na1334_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1270_1), .IN6(na679_2), .IN7(na647_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1334_2 ( .OUT(na1334_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1334_1_i) );
// C_XOR/D///      x106y98     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1335_1 ( .OUT(na1335_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na648_1), .IN6(na680_1), .IN7(na1271_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1335_2 ( .OUT(na1335_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1335_1_i) );
// C_///XOR/D      x118y87     80'hC0_EC00_80_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1336_4 ( .OUT(na1336_2_i), .IN1(na1304_1), .IN2(1'b0), .IN3(na681_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1336_5 ( .OUT(na1336_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1336_2_i) );
// C_///XOR/D      x111y65     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1337_4 ( .OUT(na1337_2_i), .IN1(na1273_1), .IN2(na650_1), .IN3(na682_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1337_5 ( .OUT(na1337_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1337_2_i) );
// C_///XOR/D      x106y65     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1338_4 ( .OUT(na1338_2_i), .IN1(~na651_2), .IN2(~na467_2), .IN3(na683_2), .IN4(na3128_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1338_5 ( .OUT(na1338_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1338_2_i) );
// C_///XOR/D      x109y76     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1339_4 ( .OUT(na1339_2_i), .IN1(na927_1), .IN2(~na468_2), .IN3(na684_1), .IN4(~na652_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1339_5 ( .OUT(na1339_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1339_2_i) );
// C_XOR/D///      x90y107     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1340_1 ( .OUT(na1340_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1244_1), .IN6(na469_2), .IN7(~na621_1),
                      .IN8(~na653_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1340_2 ( .OUT(na1340_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1340_1_i) );
// C_XOR/D///      x85y105     80'hC0_EC00_00_0000_0666_5CC9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1341_1 ( .OUT(na1341_1_i), .IN1(na654_1), .IN2(~na470_2), .IN3(1'b0), .IN4(na69_1), .IN5(1'b0), .IN6(na470_1), .IN7(~na622_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1341_2 ( .OUT(na1341_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1341_1_i) );
// C_///XOR/D      x87y94     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1342_4 ( .OUT(na1342_2_i), .IN1(~na623_1), .IN2(~na655_2), .IN3(na1246_1), .IN4(na471_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1342_5 ( .OUT(na1342_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1342_2_i) );
// C_XOR/D///      x95y78     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1343_1 ( .OUT(na1343_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na624_2), .IN6(na1247_1), .IN7(~na656_1),
                      .IN8(na472_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1343_2 ( .OUT(na1343_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1343_1_i) );
// C_///XOR/D      x92y68     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1344_4 ( .OUT(na1344_2_i), .IN1(na473_2), .IN2(na1248_1), .IN3(~na657_2), .IN4(~na625_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1344_5 ( .OUT(na1344_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1344_2_i) );
// C_XOR/D///      x101y65     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na626_2), .IN6(na1249_1), .IN7(na3032_2),
                      .IN8(~na658_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1345_2 ( .OUT(na1345_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1345_1_i) );
// C_///XOR/D      x90y66     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1346_4 ( .OUT(na1346_2_i), .IN1(na475_1), .IN2(na1250_1), .IN3(~na659_2), .IN4(~na627_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1346_5 ( .OUT(na1346_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1346_2_i) );
// C_///XOR/D      x94y67     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1347_4 ( .OUT(na1347_2_i), .IN1(1'b0), .IN2(na660_1), .IN3(na1283_1), .IN4(na3034_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1347_5 ( .OUT(na1347_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1347_2_i) );
// C_XOR/D///      x118y95     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1348_1 ( .OUT(na1348_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na629_2), .IN6(na477_1), .IN7(na1252_1),
                      .IN8(~na661_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1348_2 ( .OUT(na1348_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1348_1_i) );
// C_XOR/D///      x110y101     80'hC0_EC00_00_0000_0666_CC6A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1349_1 ( .OUT(na1349_1_i), .IN1(na739_1), .IN2(1'b0), .IN3(~na630_1), .IN4(~na478_2), .IN5(1'b0), .IN6(na662_1), .IN7(1'b0),
                      .IN8(na478_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1349_2 ( .OUT(na1349_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1349_1_i) );
// C_///XOR/D      x122y89     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1350_4 ( .OUT(na1350_2_i), .IN1(~na631_1), .IN2(na1254_1), .IN3(na479_2), .IN4(~na663_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1350_5 ( .OUT(na1350_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1350_2_i) );
// C_XOR/D///      x118y76     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_1 ( .OUT(na1351_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3039_2), .IN6(~na664_1), .IN7(na1255_1),
                      .IN8(~na632_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1351_2 ( .OUT(na1351_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1351_1_i) );
// C_///XOR/D      x117y72     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1352_4 ( .OUT(na1352_2_i), .IN1(na481_2), .IN2(~na665_2), .IN3(~na633_2), .IN4(na1256_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1352_5 ( .OUT(na1352_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1352_2_i) );
// C_XOR/D///      x113y74     80'hC0_EC00_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_1 ( .OUT(na1353_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na666_1), .IN6(1'b0), .IN7(na1289_1), .IN8(na482_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1353_2 ( .OUT(na1353_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1353_1_i) );
// C_///XOR/D      x113y71     80'hC0_EC00_80_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1354_4 ( .OUT(na1354_2_i), .IN1(na483_2), .IN2(1'b0), .IN3(na667_2), .IN4(na1290_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1354_5 ( .OUT(na1354_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1354_2_i) );
// C_///XOR/D      x117y73     80'hC0_EC00_80_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1355_4 ( .OUT(na1355_2_i), .IN1(na668_1), .IN2(na484_2), .IN3(na1291_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1355_5 ( .OUT(na1355_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1355_2_i) );
// C_XOR/D///      x118y86     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1356_1 ( .OUT(na1356_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na669_2), .IN6(na485_1), .IN7(na1260_1),
                      .IN8(~na637_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1356_2 ( .OUT(na1356_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1356_1_i) );
// C_///XOR/D      x114y80     80'hC0_EC00_80_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1357_4 ( .OUT(na1357_2_i), .IN1(~na3060_2), .IN2(na486_1), .IN3(na1261_1), .IN4(~na638_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1357_5 ( .OUT(na1357_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1357_2_i) );
// C_///XOR/D      x106y110     80'hC0_EC00_80_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1358_4 ( .OUT(na1358_2_i), .IN1(1'b0), .IN2(na487_1), .IN3(na671_2), .IN4(na1294_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1358_5 ( .OUT(na1358_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1358_2_i) );
// C_XOR/D///      x120y99     80'hC0_EC00_00_0000_0C66_6600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_1 ( .OUT(na1359_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na640_1), .IN6(~na672_1), .IN7(na1263_1),
                      .IN8(na488_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1359_2 ( .OUT(na1359_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1359_1_i) );
// C_///XOR/D      x105y108     80'hC0_EC00_80_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1360_4 ( .OUT(na1360_2_i), .IN1(na673_2), .IN2(na1296_1), .IN3(1'b0), .IN4(na489_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1360_5 ( .OUT(na1360_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1360_2_i) );
// C_XOR/D///      x119y92     80'hC0_EC00_00_0000_0666_5096
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1361_1 ( .OUT(na1361_1_i), .IN1(na842_1), .IN2(na674_1), .IN3(na490_1), .IN4(~na642_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na490_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1361_2 ( .OUT(na1361_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1361_1_i) );
// C_///XOR/D      x114y72     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1362_4 ( .OUT(na1362_2_i), .IN1(na491_2), .IN2(na1266_1), .IN3(~na675_2), .IN4(~na643_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1362_5 ( .OUT(na1362_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1362_2_i) );
// C_XOR/D///      x110y104     80'hC0_EC00_00_0000_0666_3690
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_1 ( .OUT(na1363_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na644_1), .IN4(na492_1), .IN5(na847_1), .IN6(na676_1), .IN7(1'b0),
                      .IN8(~na492_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1363_2 ( .OUT(na1363_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1363_1_i) );
// C_XOR/D///      x87y100     80'hC0_EC00_00_0000_0666_CA6C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1_i), .IN1(1'b0), .IN2(na677_2), .IN3(~na645_2), .IN4(~na461_2), .IN5(na849_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na461_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1364_2 ( .OUT(na1364_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1364_1_i) );
// C_XOR/D///      x92y110     80'hC0_EC00_00_0000_0666_6309
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1365_1 ( .OUT(na1365_1_i), .IN1(~na646_1), .IN2(na462_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na462_2), .IN7(na678_1),
                      .IN8(na899_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1365_2 ( .OUT(na1365_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1365_1_i) );
// C_XOR/D///      x92y105     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_1 ( .OUT(na1366_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na463_2), .IN6(~na679_2), .IN7(~na647_2),
                      .IN8(na3161_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1366_2 ( .OUT(na1366_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1366_1_i) );
// C_///XOR/D      x106y95     80'hC0_EC00_80_0000_0C06_FF66
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1367_4 ( .OUT(na1367_2_i), .IN1(~na648_1), .IN2(~na680_1), .IN3(na1271_1), .IN4(na3030_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0100)) 
           _a1367_5 ( .OUT(na1367_2), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1367_2_i) );
// C_XOR/D///      x113y88     80'hC0_EC00_00_0000_0C66_A600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1368_1 ( .OUT(na1368_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1304_1), .IN6(na465_1), .IN7(na681_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1368_2 ( .OUT(na1368_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1368_1_i) );
// C_XOR/D///      x110y70     80'hC0_EC00_00_0000_0C66_9900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1369_1 ( .OUT(na1369_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na466_1), .IN6(~na650_1), .IN7(~na682_1),
                      .IN8(na3162_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1369_2 ( .OUT(na1369_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1369_1_i) );
// C_XOR/D///      x103y68     80'hC0_EC00_00_0000_0666_09A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1370_1 ( .OUT(na1370_1_i), .IN1(~na651_2), .IN2(na467_1), .IN3(na683_2), .IN4(1'b0), .IN5(na925_1), .IN6(~na467_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1370_2 ( .OUT(na1370_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1370_1_i) );
// C_XOR/D///      x107y71     80'hC0_EC00_00_0000_0666_0396
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1371_1 ( .OUT(na1371_1_i), .IN1(na927_1), .IN2(na468_1), .IN3(na684_1), .IN4(~na652_1), .IN5(1'b0), .IN6(~na468_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0011_0000)) 
           _a1371_2 ( .OUT(na1371_1), .CLK(1'b0), .EN(1'b0), .SR(na2404_1), .CINY2(na3263_3), .PINY2(~na3263_6), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1371_1_i) );
// C_XOR////      x83y84     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1372_1 ( .OUT(na1372_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na55_2), .IN6(na1373_1), .IN7(~na214_2), .IN8(na2999_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y92     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1373_1 ( .OUT(na1373_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na3002_2), .IN8(na220_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x80y109     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1374_4 ( .OUT(na1374_2), .IN1(~na1376_2), .IN2(na1373_1), .IN3(na1375_2), .IN4(~na3000_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x80y103     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1375_4 ( .OUT(na1375_2), .IN1(na55_1), .IN2(1'b0), .IN3(~na129_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x81y105     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1376_4 ( .OUT(na1376_2), .IN1(na226_2), .IN2(na1455_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y90     80'h00_0018_00_0000_0666_CA6C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1377_1 ( .OUT(na1377_1), .IN1(1'b0), .IN2(na190_2), .IN3(na184_2), .IN4(na146_1), .IN5(na226_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na146_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y77     80'h00_0018_00_0000_0666_9399
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1379_1 ( .OUT(na1379_1), .IN1(~na176_2), .IN2(na190_1), .IN3(~na129_1), .IN4(na152_2), .IN5(1'b0), .IN6(~na190_2), .IN7(~na129_2),
                      .IN8(na152_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x84y71     80'h00_0018_00_0000_0666_6569
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1381_1 ( .OUT(na1381_1), .IN1(na196_1), .IN2(~na99_2), .IN3(na129_1), .IN4(na152_2), .IN5(~na196_2), .IN6(1'b0), .IN7(na129_2),
                      .IN8(na107_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y65     80'h00_0018_00_0000_0666_909C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1383_1 ( .OUT(na1383_1), .IN1(1'b0), .IN2(na202_1), .IN3(na164_1), .IN4(~na107_1), .IN5(1'b0), .IN6(1'b0), .IN7(na164_2),
                      .IN8(~na107_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x85y66     80'h00_0018_00_0000_0666_A93C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1385_1 ( .OUT(na1385_1), .IN1(1'b0), .IN2(na208_1), .IN3(1'b0), .IN4(~na256_1), .IN5(~na3007_2), .IN6(na202_2), .IN7(na164_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x84y74     80'h00_0018_00_0000_0666_CA95
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1), .IN1(~na176_1), .IN2(1'b0), .IN3(na214_1), .IN4(~na152_2), .IN5(na123_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na256_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y86     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1389_1 ( .OUT(na1389_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na176_1), .IN6(~na3009_2), .IN7(na1375_2),
                      .IN8(na220_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x81y92     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1390_4 ( .OUT(na1390_2), .IN1(na1376_2), .IN2(~na1391_2), .IN3(na1375_2), .IN4(~na146_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x83y84     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1391_4 ( .OUT(na1391_2), .IN1(na55_2), .IN2(1'b0), .IN3(~na3004_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y85     80'h00_0018_00_0000_0666_AA39
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1392_1 ( .OUT(na1392_1), .IN1(na140_1), .IN2(~na190_2), .IN3(1'b0), .IN4(~na146_2), .IN5(na176_2), .IN6(1'b0), .IN7(na184_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x84y79     80'h00_0018_00_0000_0666_A996
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1394_1 ( .OUT(na1394_1), .IN1(na176_1), .IN2(na99_2), .IN3(na129_2), .IN4(~na146_1), .IN5(~na176_2), .IN6(na190_1), .IN7(na129_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y72     80'h00_0018_00_0000_0666_9A69
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1396_1 ( .OUT(na1396_1), .IN1(na196_1), .IN2(~na99_2), .IN3(na129_1), .IN4(na152_1), .IN5(na176_1), .IN6(1'b0), .IN7(~na2995_2),
                      .IN8(na107_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x84y68     80'h00_0018_00_0000_0666_0693
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1398_1 ( .OUT(na1398_1), .IN1(1'b0), .IN2(~na202_2), .IN3(~na164_2), .IN4(na107_1), .IN5(na196_2), .IN6(na202_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y65     80'h00_0018_00_0000_0666_ACC6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1400_1 ( .OUT(na1400_1), .IN1(na123_1), .IN2(na202_2), .IN3(1'b0), .IN4(na256_1), .IN5(1'b0), .IN6(na208_1), .IN7(na164_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y72     80'h00_0018_00_0000_0666_A59C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1402_1 ( .OUT(na1402_1), .IN1(1'b0), .IN2(na208_2), .IN3(na129_1), .IN4(~na152_2), .IN5(~na123_1), .IN6(1'b0), .IN7(na214_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y86     80'h00_0018_00_0000_0C66_9600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1404_1 ( .OUT(na1404_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na55_1), .IN6(na1391_2), .IN7(na214_1), .IN8(~na220_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y87     80'h00_0018_00_0000_0666_66A5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1405_1 ( .OUT(na1405_1), .IN1(~na140_1), .IN2(1'b0), .IN3(na214_1), .IN4(1'b0), .IN5(na226_2), .IN6(na1391_2), .IN7(na214_2),
                      .IN8(na146_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x80y90     80'h00_0018_00_0000_0666_C909
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1407_1 ( .OUT(na1407_1), .IN1(~na140_1), .IN2(na1455_1), .IN3(1'b0), .IN4(1'b0), .IN5(na176_2), .IN6(~na190_2), .IN7(1'b0),
                      .IN8(na146_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y81     80'h00_0018_00_0000_0666_969A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1409_1 ( .OUT(na1409_1), .IN1(na176_1), .IN2(1'b0), .IN3(na129_2), .IN4(~na146_1), .IN5(na3008_2), .IN6(na99_2), .IN7(na184_2),
                      .IN8(~na152_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y78     80'h00_0018_00_0000_0666_6963
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_1 ( .OUT(na1411_1), .IN1(1'b0), .IN2(~na190_1), .IN3(na214_1), .IN4(na107_1), .IN5(~na196_2), .IN6(na3001_2), .IN7(na3003_2),
                      .IN8(na107_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y69     80'h00_0018_00_0000_0666_A5A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1413_1 ( .OUT(na1413_1), .IN1(na196_1), .IN2(~na202_2), .IN3(na164_2), .IN4(1'b0), .IN5(~na196_2), .IN6(1'b0), .IN7(na164_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x85y67     80'h00_0018_00_0000_0666_C95C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1414_1 ( .OUT(na1414_1), .IN1(1'b0), .IN2(na202_1), .IN3(~na164_1), .IN4(1'b0), .IN5(na123_1), .IN6(~na208_2), .IN7(1'b0),
                      .IN8(na256_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y74     80'h00_0018_00_0000_0666_9306
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1415_1 ( .OUT(na1415_1), .IN1(na176_1), .IN2(na208_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na208_2), .IN7(~na129_1),
                      .IN8(na152_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y83     80'h00_0018_00_0000_0666_AA95
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1417_1 ( .OUT(na1417_1), .IN1(~na55_2), .IN2(1'b0), .IN3(~na214_2), .IN4(na152_2), .IN5(na55_1), .IN6(1'b0), .IN7(na214_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y94     80'h00_0018_00_0000_0666_6CA9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1419_1 ( .OUT(na1419_1), .IN1(na140_1), .IN2(~na1455_1), .IN3(na214_1), .IN4(1'b0), .IN5(1'b0), .IN6(na1373_1), .IN7(na214_2),
                      .IN8(na146_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x81y89     80'h00_0060_00_0000_0C06_FF99
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1420_4 ( .OUT(na1420_2), .IN1(na1376_2), .IN2(~na3005_2), .IN3(na184_2), .IN4(~na146_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y80     80'h00_0018_00_0000_0666_969C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1421_1 ( .OUT(na1421_1), .IN1(1'b0), .IN2(na190_2), .IN3(na184_2), .IN4(~na152_2), .IN5(na2991_2), .IN6(na190_1), .IN7(na214_1),
                      .IN8(~na152_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x84y75     80'h00_0018_00_0000_0666_6A66
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1423_1 ( .OUT(na1423_1), .IN1(~na196_1), .IN2(~na190_1), .IN3(na214_1), .IN4(na107_1), .IN5(na196_2), .IN6(1'b0), .IN7(na129_2),
                      .IN8(na152_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y68     80'h00_0018_00_0000_0666_0963
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1425_1 ( .OUT(na1425_1), .IN1(1'b0), .IN2(~na202_1), .IN3(na164_1), .IN4(na107_2), .IN5(na196_1), .IN6(~na202_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x86y67     80'h00_0018_00_0000_0666_C3A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1427_1 ( .OUT(na1427_1), .IN1(na123_1), .IN2(~na208_1), .IN3(na164_2), .IN4(1'b0), .IN5(1'b0), .IN6(~na208_2), .IN7(1'b0),
                      .IN8(na3006_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x84y73     80'h00_0018_00_0000_0666_A099
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1428_1 ( .OUT(na1428_1), .IN1(~na176_1), .IN2(na208_1), .IN3(na129_1), .IN4(~na256_1), .IN5(1'b0), .IN6(1'b0), .IN7(na214_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y104     80'h00_0018_00_0040_0AE9_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1436_1 ( .OUT(na1436_1), .IN1(na3170_2), .IN2(1'b1), .IN3(~na2409_2), .IN4(1'b1), .IN5(1'b1), .IN6(na2413_2), .IN7(na2409_1),
                      .IN8(~na2964_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x80y100     80'h00_0018_00_0040_0C49_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1438_1 ( .OUT(na1438_1), .IN1(na2930_1), .IN2(1'b0), .IN3(1'b1), .IN4(na3218_2), .IN5(1'b1), .IN6(~na1023_1), .IN7(1'b1),
                      .IN8(na1029_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x80y103     80'h00_0018_00_0000_0C66_3D00
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1439_1 ( .OUT(na1439_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2931_2), .IN6(~na23_2), .IN7(1'b1), .IN8(na1021_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y108     80'h00_0018_00_0040_0AB0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1440_1 ( .OUT(na1440_1), .IN1(1'b1), .IN2(na23_1), .IN3(1'b1), .IN4(na2410_2), .IN5(na20_2), .IN6(na2933_1), .IN7(1'b0),
                      .IN8(na25_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y93     80'h00_0018_00_0000_0666_A069
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1443_1 ( .OUT(na1443_1), .IN1(na18_1), .IN2(~na23_2), .IN3(~na2934_2), .IN4(~na32_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2934_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y75     80'h00_0018_00_0040_0AE5_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1444_1 ( .OUT(na1444_1), .IN1(1'b1), .IN2(~na2428_2), .IN3(na1018_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2428_1), .IN7(~na36_1),
                      .IN8(na35_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y97     80'h00_0018_00_0040_0A3F_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1446_1 ( .OUT(na1446_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(~na1656_2), .IN6(~na819_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x100y93     80'h00_0018_00_0040_0A3F_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1448_1 ( .OUT(na1448_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(~na2236_2), .IN6(~na961_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y93     80'h00_0018_00_0000_0EEE_DC53
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1449_1 ( .OUT(na1449_1), .IN1(1'b0), .IN2(~na2936_2), .IN3(~na1446_1), .IN4(1'b0), .IN5(1'b0), .IN6(na182_1), .IN7(~na1448_1),
                      .IN8(na2937_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x105y94     80'h00_0018_00_0040_0A3F_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1), .IN1(na1087_2), .IN2(1'b1), .IN3(na1103_2), .IN4(1'b1), .IN5(~na1657_1), .IN6(~na828_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y89     80'h00_0018_00_0040_0A3F_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1453_1 ( .OUT(na1453_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2982_2), .IN5(~na962_1), .IN6(~na2237_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x98y93     80'h00_0018_00_0000_0EEE_C55B
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1454_1 ( .OUT(na1454_1), .IN1(na183_1), .IN2(~na1451_1), .IN3(~na2939_2), .IN4(1'b0), .IN5(~na1453_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na2940_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x85y92     80'h40_E800_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1455_1 ( .OUT(na1455_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1454_1), .IN8(~na2986_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1455_2 ( .OUT(na1455_1), .CLK(1'b0), .EN(na429_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1455_1_i) );
// C_XOR////      x124y86     80'h00_0018_00_0000_0C66_C300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1456_1 ( .OUT(na1456_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na707_1), .IN7(1'b0), .IN8(na2942_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x123y79     80'h00_0060_00_0000_0C06_FF3E
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1457_4 ( .OUT(na1457_2), .IN1(~na3074_2), .IN2(~na704_1), .IN3(1'b1), .IN4(na1456_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x125y75     80'h00_0018_00_0000_0C66_EAFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1458_1 ( .OUT(na1458_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1457_2), .IN6(1'b1), .IN7(~na706_1), .IN8(~na702_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y101     80'h00_0018_00_0040_0AFC_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1459_1 ( .OUT(na1459_1), .IN1(1'b1), .IN2(~na3096_2), .IN3(1'b1), .IN4(na784_1), .IN5(na3095_2), .IN6(na779_1), .IN7(~na780_2),
                      .IN8(~na3094_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x121y100     80'h00_0060_00_0000_0C06_FF5E
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1460_4 ( .OUT(na1460_2), .IN1(~na3098_2), .IN2(~na2716_2), .IN3(na1459_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x124y100     80'h00_0018_00_0000_0C66_ECFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1461_1 ( .OUT(na1461_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1460_2), .IN7(~na783_1), .IN8(~na781_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y89     80'h00_0018_00_0040_0A7A_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1462_1 ( .OUT(na1462_1), .IN1(1'b1), .IN2(~na2716_2), .IN3(1'b1), .IN4(na2722_2), .IN5(na3141_2), .IN6(~na2716_1), .IN7(na780_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x116y112     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1464_1 ( .OUT(na1464_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na858_2), .IN5(na856_1), .IN6(1'b0), .IN7(na2950_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y109     80'h00_0018_00_0000_0666_A365
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1465_1 ( .OUT(na1465_1), .IN1(~na3201_2), .IN2(1'b0), .IN3(na2748_2), .IN4(na1464_1), .IN5(1'b0), .IN6(~na862_1), .IN7(na2748_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x113y105     80'h00_0018_00_0040_0A78_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1466_1 ( .OUT(na1466_1), .IN1(1'b1), .IN2(~na1067_1), .IN3(na2769_2), .IN4(1'b1), .IN5(na853_1), .IN6(na2951_1), .IN7(na877_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x117y99     80'h00_0018_00_0000_0666_FDB5
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1467_1 ( .OUT(na1467_1), .IN1(na1466_1), .IN2(1'b1), .IN3(~na878_1), .IN4(na882_1), .IN5(na3121_2), .IN6(~na883_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y86     80'h00_0078_00_0020_0C66_3530
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1469_1 ( .OUT(na1469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na2961_2),
                      .CINX(1'b0), .CINY1(na1474_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1469_4 ( .OUT(na1469_2), .COUTY1(na1469_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na7_1), .IN5(~na6_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na2961_2), .CINX(1'b0), .CINY1(na1474_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y87     80'h00_0078_00_0020_0C66_5005
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1471_1 ( .OUT(na1471_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1469_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1471_4 ( .OUT(na1471_2), .COUTY1(na1471_4), .IN1(~na6_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na8_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1469_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y88     80'h00_0018_00_0010_0666_0003
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1473_1 ( .OUT(na1473_1), .COUTY1(na1473_4), .IN1(1'b1), .IN2(~na5_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na1471_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x93y85     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1474_2 ( .OUT(na1474_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1474_6 ( .COUTY1(na1474_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1474_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x97y79     80'h00_0078_00_0020_0C66_CC0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1475_1 ( .OUT(na1475_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na5_1), .IN7(1'b1), .IN8(na7_2),
                      .CINX(1'b0), .CINY1(na1481_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1475_4 ( .OUT(na1475_2), .COUTY1(na1475_4), .IN1(na6_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na5_1), .IN7(1'b1),
                      .IN8(na7_2), .CINX(1'b0), .CINY1(na1481_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y80     80'h00_0078_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1477_1 ( .OUT(na1477_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na7_1),
                      .CINX(1'b0), .CINY1(na1475_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1477_4 ( .OUT(na1477_2), .COUTY1(na1477_4), .IN1(1'b0), .IN2(1'b0), .IN3(na8_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na7_1), .CINX(1'b0), .CINY1(na1475_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y81     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1479_1 ( .OUT(na1479_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na6_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1477_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1479_4 ( .OUT(na1479_2), .IN1(1'b1), .IN2(na5_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1477_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x97y78     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1481_2 ( .OUT(na1481_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1481_6 ( .COUTY1(na1481_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1481_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x110y95     80'h00_0078_00_0020_0C66_AAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1482_1 ( .OUT(na1482_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1087_2), .IN6(1'b1), .IN7(na1089_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na2411_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1482_4 ( .OUT(na1482_2), .COUTY1(na1482_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1089_1), .IN4(1'b1), .IN5(na1087_2), .IN6(1'b1),
                      .IN7(na1089_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na2411_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x110y96     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1484_1 ( .OUT(na1484_1), .IN1(1'b1), .IN2(na1090_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1482_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0018_0018)) 
           _a1487 ( .GLB0(na1487_1), .GLB1(na1487_2), .GLB2(_d0), .GLB3(_d1), .CLK_FB0(_d2), .CLK_FB1(_d3), .CLK_FB2(_d4), .CLK_FB3(_d5),
                    .CLK0_0(1'b0), .CLK0_90(1'b0), .CLK0_180(1'b0), .CLK0_270(1'b0), .CLK0_BYP(1'b0), .CLK1_0(1'b0), .CLK1_90(1'b0),
                    .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                    .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(na1489_9),
                    .USR_GLB1(na1488_9), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_AND////      x1y127     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1488_1 ( .OUT(na1488_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2395_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1488_6 ( .RAM_O1(na1488_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1488_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x1y128     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1489_1 ( .OUT(na1489_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1114_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1489_6 ( .RAM_O1(na1489_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1489_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/D      x86y92     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1592_4 ( .OUT(na1592_2_i), .IN1(na1009_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1592_5 ( .OUT(na1592_2), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1592_2_i) );
// C_AND/D///      x83y101     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1593_1 ( .OUT(na1593_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1011_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1593_2 ( .OUT(na1593_1), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1593_1_i) );
// C_///AND/D      x87y92     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1594_4 ( .OUT(na1594_2_i), .IN1(na1012_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1594_5 ( .OUT(na1594_2), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1594_2_i) );
// C_AND/D///      x90y85     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1595_1 ( .OUT(na1595_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1013_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1595_2 ( .OUT(na1595_1), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1595_1_i) );
// C_///AND/D      x87y82     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1596_4 ( .OUT(na1596_2_i), .IN1(na1014_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1596_5 ( .OUT(na1596_2), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1596_2_i) );
// C_AND/D///      x89y71     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1597_1 ( .OUT(na1597_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1015_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1597_2 ( .OUT(na1597_1), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1597_1_i) );
// C_///AND/D      x91y78     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1598_4 ( .OUT(na1598_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1016_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1598_5 ( .OUT(na1598_2), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1598_2_i) );
// C_AND/D///      x90y76     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_1 ( .OUT(na1599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1017_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1599_2 ( .OUT(na1599_1), .CLK(1'b0), .EN(na82_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1599_1_i) );
// C_///AND/D      x117y81     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1624_4 ( .OUT(na1624_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na693_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1624_5 ( .OUT(na1624_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1624_2_i) );
// C_AND/D///      x105y95     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1625_1 ( .OUT(na1625_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na739_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1625_2 ( .OUT(na1625_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1625_1_i) );
// C_///AND/D      x107y89     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1626_4 ( .OUT(na1626_2_i), .IN1(na748_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1626_5 ( .OUT(na1626_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1626_2_i) );
// C_AND/D///      x105y77     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1627_1 ( .OUT(na1627_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na754_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1627_2 ( .OUT(na1627_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1627_1_i) );
// C_///AND/D      x98y79     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1628_4 ( .OUT(na1628_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na760_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1628_5 ( .OUT(na1628_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1628_2_i) );
// C_AND/D///      x102y65     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1629_1 ( .OUT(na1629_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na764_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1629_2 ( .OUT(na1629_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1629_1_i) );
// C_///AND/D      x99y67     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1630_4 ( .OUT(na1630_2_i), .IN1(na769_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1630_5 ( .OUT(na1630_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1630_2_i) );
// C_AND/D///      x99y67     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1631_1 ( .OUT(na1631_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na771_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1631_2 ( .OUT(na1631_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1631_1_i) );
// C_///AND/D      x93y104     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1640_4 ( .OUT(na1640_2_i), .IN1(na849_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1640_5 ( .OUT(na1640_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1640_2_i) );
// C_AND/D///      x96y110     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1641_1 ( .OUT(na1641_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na899_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1641_2 ( .OUT(na1641_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1641_1_i) );
// C_///AND/D      x99y101     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1642_4 ( .OUT(na1642_2_i), .IN1(1'b1), .IN2(na908_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1642_5 ( .OUT(na1642_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1642_2_i) );
// C_AND/D///      x97y94     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1643_1 ( .OUT(na1643_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na912_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1643_2 ( .OUT(na1643_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1643_1_i) );
// C_///AND/D      x96y93     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1644_4 ( .OUT(na1644_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na918_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1644_5 ( .OUT(na1644_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1644_2_i) );
// C_AND/D///      x110y84     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1645_1 ( .OUT(na1645_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na921_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1645_2 ( .OUT(na1645_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1645_1_i) );
// C_///AND/D      x104y78     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1646_4 ( .OUT(na1646_2_i), .IN1(na925_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1646_5 ( .OUT(na1646_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1646_2_i) );
// C_AND/D///      x105y82     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1647_1 ( .OUT(na1647_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na927_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1647_2 ( .OUT(na1647_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1647_1_i) );
// C_///AND/D      x107y99     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1648_4 ( .OUT(na1648_2_i), .IN1(1'b1), .IN2(na774_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1648_5 ( .OUT(na1648_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1648_2_i) );
// C_AND/D///      x108y93     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1649_1 ( .OUT(na1649_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na820_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1649_2 ( .OUT(na1649_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1649_1_i) );
// C_///AND/D      x91y110     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1650_4 ( .OUT(na1650_2_i), .IN1(na829_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1650_5 ( .OUT(na1650_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1650_2_i) );
// C_AND/D///      x89y103     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1651_1 ( .OUT(na1651_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na833_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1651_2 ( .OUT(na1651_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1651_1_i) );
// C_///AND/D      x99y107     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1652_4 ( .OUT(na1652_2_i), .IN1(na839_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1652_5 ( .OUT(na1652_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1652_2_i) );
// C_AND/D///      x115y95     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1653_1 ( .OUT(na1653_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na842_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1653_2 ( .OUT(na1653_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1653_1_i) );
// C_///AND/D      x113y89     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1654_4 ( .OUT(na1654_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na845_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1654_5 ( .OUT(na1654_2), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1654_2_i) );
// C_AND/D///      x106y105     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1655_1 ( .OUT(na1655_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na847_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1655_2 ( .OUT(na1655_1), .CLK(1'b0), .EN(na65_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1655_1_i) );
// C_///AND/D      x107y97     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1656_4 ( .OUT(na1656_2_i), .IN1(1'b1), .IN2(na774_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1656_5 ( .OUT(na1656_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1656_2_i) );
// C_AND/D///      x113y95     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1657_1 ( .OUT(na1657_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na820_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1657_2 ( .OUT(na1657_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1657_1_i) );
// C_///AND/D      x90y111     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1658_4 ( .OUT(na1658_2_i), .IN1(na829_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1658_5 ( .OUT(na1658_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1658_2_i) );
// C_AND/D///      x89y104     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1659_1 ( .OUT(na1659_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na833_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1659_2 ( .OUT(na1659_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1659_1_i) );
// C_///AND/D      x98y105     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1660_4 ( .OUT(na1660_2_i), .IN1(na839_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1660_5 ( .OUT(na1660_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1660_2_i) );
// C_AND/D///      x116y95     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1661_1 ( .OUT(na1661_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na842_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1661_2 ( .OUT(na1661_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1661_1_i) );
// C_///AND/D      x111y91     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1662_4 ( .OUT(na1662_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na845_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1662_5 ( .OUT(na1662_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1662_2_i) );
// C_AND/D///      x105y104     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1663_1 ( .OUT(na1663_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na847_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1663_2 ( .OUT(na1663_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1663_1_i) );
// C_///AND/D      x116y84     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1664_4 ( .OUT(na1664_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na693_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1664_5 ( .OUT(na1664_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1664_2_i) );
// C_AND/D///      x106y96     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1665_1 ( .OUT(na1665_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na739_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1665_2 ( .OUT(na1665_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1665_1_i) );
// C_///AND/D      x104y86     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1666_4 ( .OUT(na1666_2_i), .IN1(na748_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1666_5 ( .OUT(na1666_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1666_2_i) );
// C_AND/D///      x104y76     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1667_1 ( .OUT(na1667_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na754_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1667_2 ( .OUT(na1667_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1667_1_i) );
// C_///AND/D      x100y72     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1668_4 ( .OUT(na1668_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na760_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1668_5 ( .OUT(na1668_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1668_2_i) );
// C_AND/D///      x103y64     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1669_1 ( .OUT(na1669_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na764_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1669_2 ( .OUT(na1669_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1669_1_i) );
// C_///AND/D      x97y66     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1670_4 ( .OUT(na1670_2_i), .IN1(na769_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1670_5 ( .OUT(na1670_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1670_2_i) );
// C_AND/D///      x102y67     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1671_1 ( .OUT(na1671_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na771_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1671_2 ( .OUT(na1671_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1671_1_i) );
// C_///AND/D      x84y101     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1672_4 ( .OUT(na1672_2_i), .IN1(na11_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1672_5 ( .OUT(na1672_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1672_2_i) );
// C_AND/D///      x81y102     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1673_1 ( .OUT(na1673_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na69_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1673_2 ( .OUT(na1673_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1673_1_i) );
// C_///AND/D      x85y85     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1674_4 ( .OUT(na1674_2_i), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1674_5 ( .OUT(na1674_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1674_2_i) );
// C_AND/D///      x85y81     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1675_1 ( .OUT(na1675_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na94_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1675_2 ( .OUT(na1675_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1675_1_i) );
// C_///AND/D      x89y79     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1676_4 ( .OUT(na1676_2_i), .IN1(1'b1), .IN2(na105_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1676_5 ( .OUT(na1676_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1676_2_i) );
// C_AND/D///      x91y70     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1677_1 ( .OUT(na1677_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na112_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1677_2 ( .OUT(na1677_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1677_1_i) );
// C_///AND/D      x89y75     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1678_4 ( .OUT(na1678_2_i), .IN1(na121_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1678_5 ( .OUT(na1678_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1678_2_i) );
// C_AND/D///      x87y72     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1679_1 ( .OUT(na1679_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na128_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1679_2 ( .OUT(na1679_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1679_1_i) );
// C_///AND/D      x84y102     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1680_4 ( .OUT(na1680_2_i), .IN1(na849_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1680_5 ( .OUT(na1680_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1680_2_i) );
// C_AND/D///      x91y108     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1681_1 ( .OUT(na1681_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na899_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1681_2 ( .OUT(na1681_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1681_1_i) );
// C_///AND/D      x97y104     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1682_4 ( .OUT(na1682_2_i), .IN1(1'b1), .IN2(na908_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1682_5 ( .OUT(na1682_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1682_2_i) );
// C_AND/D///      x93y93     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1683_1 ( .OUT(na1683_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na912_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1683_2 ( .OUT(na1683_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1683_1_i) );
// C_///AND/D      x93y90     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1684_4 ( .OUT(na1684_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na918_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1684_5 ( .OUT(na1684_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1684_2_i) );
// C_AND/D///      x101y88     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1685_1 ( .OUT(na1685_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na921_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1685_2 ( .OUT(na1685_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1685_1_i) );
// C_///AND/D      x98y71     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1686_4 ( .OUT(na1686_2_i), .IN1(na925_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a1686_5 ( .OUT(na1686_2), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1686_2_i) );
// C_AND/D///      x101y81     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1687_1 ( .OUT(na1687_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na927_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a1687_2 ( .OUT(na1687_1), .CLK(1'b0), .EN(na82_1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1687_1_i) );
// C_///AND/D      x83y104     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2220_4 ( .OUT(na2220_2_i), .IN1(na11_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2220_5 ( .OUT(na2220_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2220_2_i) );
// C_AND/D///      x81y103     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2221_1 ( .OUT(na2221_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na69_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2221_2 ( .OUT(na2221_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2221_1_i) );
// C_///AND/D      x85y87     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2222_4 ( .OUT(na2222_2_i), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2222_5 ( .OUT(na2222_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2222_2_i) );
// C_AND/D///      x83y82     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2223_1 ( .OUT(na2223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na94_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2223_2 ( .OUT(na2223_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2223_1_i) );
// C_///AND/D      x86y75     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2224_4 ( .OUT(na2224_2_i), .IN1(1'b1), .IN2(na105_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2224_5 ( .OUT(na2224_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2224_2_i) );
// C_AND/D///      x89y69     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2225_1 ( .OUT(na2225_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na112_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2225_2 ( .OUT(na2225_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2225_1_i) );
// C_///AND/D      x88y73     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2226_4 ( .OUT(na2226_2_i), .IN1(na121_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2226_5 ( .OUT(na2226_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2226_2_i) );
// C_AND/D///      x85y72     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2227_1 ( .OUT(na2227_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na128_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2227_2 ( .OUT(na2227_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2227_1_i) );
// C_///AND/D      x84y103     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2228_4 ( .OUT(na2228_2_i), .IN1(na849_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2228_5 ( .OUT(na2228_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2228_2_i) );
// C_AND/D///      x95y108     80'h40_E800_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2229_1 ( .OUT(na2229_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na899_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2229_2 ( .OUT(na2229_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2229_1_i) );
// C_///AND/D      x95y108     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2230_4 ( .OUT(na2230_2_i), .IN1(1'b1), .IN2(na908_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2230_5 ( .OUT(na2230_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2230_2_i) );
// C_AND/D///      x93y95     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2231_1 ( .OUT(na2231_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na912_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2231_2 ( .OUT(na2231_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2231_1_i) );
// C_///AND/D      x96y94     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2232_4 ( .OUT(na2232_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na918_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2232_5 ( .OUT(na2232_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2232_2_i) );
// C_AND/D///      x105y84     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2233_1 ( .OUT(na2233_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na921_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2233_2 ( .OUT(na2233_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2233_1_i) );
// C_///AND/D      x98y65     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2234_4 ( .OUT(na2234_2_i), .IN1(na925_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2234_5 ( .OUT(na2234_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2234_2_i) );
// C_AND/D///      x100y81     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2235_1 ( .OUT(na2235_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na927_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2235_2 ( .OUT(na2235_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2235_1_i) );
// C_///AND/D      x109y97     80'h40_E800_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2236_4 ( .OUT(na2236_2_i), .IN1(1'b1), .IN2(na774_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2236_5 ( .OUT(na2236_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2236_2_i) );
// C_AND/D///      x117y100     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2237_1 ( .OUT(na2237_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na820_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2237_2 ( .OUT(na2237_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2237_1_i) );
// C_///AND/D      x91y109     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2238_4 ( .OUT(na2238_2_i), .IN1(na829_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2238_5 ( .OUT(na2238_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2238_2_i) );
// C_AND/D///      x96y101     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2239_1 ( .OUT(na2239_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na833_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2239_2 ( .OUT(na2239_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2239_1_i) );
// C_///AND/D      x96y105     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2240_4 ( .OUT(na2240_2_i), .IN1(na839_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2240_5 ( .OUT(na2240_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2240_2_i) );
// C_AND/D///      x117y95     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2241_1 ( .OUT(na2241_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na842_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2241_2 ( .OUT(na2241_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2241_1_i) );
// C_///AND/D      x117y89     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2242_4 ( .OUT(na2242_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na845_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2242_5 ( .OUT(na2242_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2242_2_i) );
// C_AND/D///      x109y103     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2243_1 ( .OUT(na2243_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na847_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2243_2 ( .OUT(na2243_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2243_1_i) );
// C_///AND/D      x117y82     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2244_4 ( .OUT(na2244_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na693_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2244_5 ( .OUT(na2244_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2244_2_i) );
// C_AND/D///      x109y89     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2245_1 ( .OUT(na2245_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na739_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2245_2 ( .OUT(na2245_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2245_1_i) );
// C_///AND/D      x105y83     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2246_4 ( .OUT(na2246_2_i), .IN1(na748_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2246_5 ( .OUT(na2246_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2246_2_i) );
// C_AND/D///      x103y75     80'h40_E800_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2247_1 ( .OUT(na2247_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na754_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2247_2 ( .OUT(na2247_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2247_1_i) );
// C_///AND/D      x98y77     80'h40_E800_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2248_4 ( .OUT(na2248_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na760_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2248_5 ( .OUT(na2248_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2248_2_i) );
// C_AND/D///      x105y65     80'h40_E800_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2249_1 ( .OUT(na2249_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na764_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2249_2 ( .OUT(na2249_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2249_1_i) );
// C_///AND/D      x97y69     80'h40_E800_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2250_4 ( .OUT(na2250_2_i), .IN1(na769_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2250_5 ( .OUT(na2250_2), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2250_2_i) );
// C_AND/D///      x102y69     80'h40_E800_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2251_1 ( .OUT(na2251_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na771_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2251_2 ( .OUT(na2251_1), .CLK(1'b0), .EN(na1010_2), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2251_1_i) );
// C_///AND/D      x89y84     80'h40_EC00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2348_4 ( .OUT(na2348_2_i), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2348_5 ( .OUT(na2348_2), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2348_2_i) );
// C_AND/D///      x89y84     80'h40_EC00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2349_1 ( .OUT(na2349_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1089_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2349_2 ( .OUT(na2349_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2349_1_i) );
// C_///AND/D      x88y84     80'h40_EC00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2350_4 ( .OUT(na2350_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1089_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0100)) 
           _a2350_5 ( .OUT(na2350_2), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2350_2_i) );
// C_AND/D///      x88y83     80'h40_EC00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2351_1 ( .OUT(na2351_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1090_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0001_0000)) 
           _a2351_2 ( .OUT(na2351_1), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2351_1_i) );
// C_MX2b////      x88y87     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2363_1 ( .OUT(na2363_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na55_1), .IN6(na1372_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x82y96     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2364_1 ( .OUT(na2364_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1374_2), .IN8(na146_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y85     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2365_1 ( .OUT(na2365_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na176_2), .IN6(na1377_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y82     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2366_1 ( .OUT(na2366_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1379_1), .IN6(na99_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y76     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2367_1 ( .OUT(na2367_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1381_1), .IN8(na107_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y70     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2368_1 ( .OUT(na2368_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1383_1), .IN6(na202_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2369_1 ( .OUT(na2369_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na123_1), .IN6(na1385_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y76     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2370_1 ( .OUT(na2370_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na129_1), .IN8(na1387_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y86     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2371_1 ( .OUT(na2371_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na55_2), .IN6(na1389_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y90     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2372_1 ( .OUT(na2372_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na140_1), .IN6(na1390_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y85     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2373_1 ( .OUT(na2373_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1392_1), .IN8(na146_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y78     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2374_1 ( .OUT(na2374_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1394_1), .IN8(na152_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y74     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2375_1 ( .OUT(na2375_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na196_2), .IN6(na1396_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y70     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2376_1 ( .OUT(na2376_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na164_1), .IN8(na1398_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y69     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2377_1 ( .OUT(na2377_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1400_1), .IN6(na208_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y73     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2378_1 ( .OUT(na2378_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na176_1), .IN6(na1402_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y86     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2379_1 ( .OUT(na2379_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na214_2), .IN8(na1404_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y83     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2380_1 ( .OUT(na2380_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1405_1), .IN6(na1455_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y95     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2381_1 ( .OUT(na2381_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na184_2), .IN8(na1407_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y89     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2382_1 ( .OUT(na2382_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1409_1), .IN6(na190_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x86y84     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2383_1 ( .OUT(na2383_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na196_1), .IN6(na1411_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y73     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2384_1 ( .OUT(na2384_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1413_1), .IN6(na202_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y73     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2385_1 ( .OUT(na2385_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1414_1), .IN6(na208_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y88     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2386_1 ( .OUT(na2386_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na214_1), .IN8(na1415_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y86     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2387_1 ( .OUT(na2387_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1417_1), .IN8(na220_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y96     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2388_1 ( .OUT(na2388_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na226_2), .IN6(na1419_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y93     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2389_1 ( .OUT(na2389_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1420_2), .IN6(na190_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y82     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2390_1 ( .OUT(na2390_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na129_2), .IN8(na1421_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y79     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2391_1 ( .OUT(na2391_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1423_1), .IN8(na107_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y72     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2392_1 ( .OUT(na2392_1), .IN1(1'b1), .IN2(na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na164_2), .IN8(na1425_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y70     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2393_1 ( .OUT(na2393_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1427_1), .IN8(na256_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x86y78     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2394_1 ( .OUT(na2394_1), .IN1(1'b1), .IN2(~na1113_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1428_1), .IN8(na152_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2395 ( .Y(na2395_1), .I(clk10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2396 ( .O(led[0]), .A(na2952_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2397 ( .O(led[1]), .A(na2953_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2398 ( .O(led[2]), .A(na2954_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2399 ( .O(led[3]), .A(na2955_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2400 ( .O(led[4]), .A(na2956_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2401 ( .O(led[5]), .A(na2957_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2402 ( .O(led[6]), .A(na2958_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a2403 ( .O(led[7]), .A(na2959_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a2404 ( .Y(na2404_1), .I(reset_n) );
// C_AND///AND/      x81y79     80'h00_0078_00_0000_0C88_CC53
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2405_1 ( .OUT(na2405_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na15_1), .IN7(1'b1), .IN8(na2967_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2405_4 ( .OUT(na2405_2), .IN1(1'b1), .IN2(~na23_2), .IN3(~na33_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x80y88     80'h00_0078_00_0000_0C66_096C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2407_1 ( .OUT(na2407_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na27_1), .IN6(na2414_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2407_4 ( .OUT(na2407_2), .IN1(1'b0), .IN2(na1440_1), .IN3(na1439_1), .IN4(na1438_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/DST      x83y110     80'h60_BC00_80_0000_0C08_FF00
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2408_4 ( .OUT(na2408_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0101_0100)) 
           _a2408_5 ( .OUT(na2408_2), .CLK(1'b0), .EN(1'b1), .SR(na2404_1), .CINY2(na3263_3), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2408_2_i) );
// C_XOR///XOR/      x80y97     80'h00_0078_00_0000_0C66_063A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2409_1 ( .OUT(na2409_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na18_1), .IN6(na2413_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2409_4 ( .OUT(na2409_2), .IN1(na1033_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1029_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x82y102     80'h00_0078_00_0000_0C66_AA63
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2410_1 ( .OUT(na2410_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na20_1), .IN6(1'b0), .IN7(na2966_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2410_4 ( .OUT(na2410_2), .IN1(1'b0), .IN2(~na1031_1), .IN3(na1027_1), .IN4(na1029_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x110y94     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a2411_2 ( .OUT(na2411_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a2411_6 ( .COUTY1(na2411_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na2411_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x93y89     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a2412_1 ( .OUT(na2412_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1473_4), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x79y100     80'h00_0078_00_0000_0C66_5CA3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2413_1 ( .OUT(na2413_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na23_2), .IN7(~na1018_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2413_4 ( .OUT(na2413_2), .IN1(1'b0), .IN2(~na1023_1), .IN3(na1027_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x79y90     80'h00_0078_00_0000_0C66_35C6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2414_1 ( .OUT(na2414_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na27_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na2407_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2414_4 ( .OUT(na2414_2), .IN1(na19_1), .IN2(na1436_1), .IN3(1'b0), .IN4(na22_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x80y70     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2416_4 ( .OUT(na2416_2), .IN1(na1443_1), .IN2(na2414_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y88     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2418_1 ( .OUT(na2418_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1443_1), .IN6(1'b0), .IN7(1'b0), .IN8(na2407_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x79y75     80'h00_0078_00_0000_0C66_A5C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2423_1 ( .OUT(na2423_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na42_2), .IN6(1'b0), .IN7(na36_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2423_4 ( .OUT(na2423_2), .IN1(~na48_1), .IN2(1'b0), .IN3(1'b0), .IN4(na25_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x77y87     80'h00_0060_00_0000_0C06_FFA3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2425_4 ( .OUT(na2425_2), .IN1(1'b0), .IN2(~na23_1), .IN3(na36_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x80y96     80'h00_0078_00_0000_0C88_F85A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2426_1 ( .OUT(na2426_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na48_2), .IN6(na15_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2426_4 ( .OUT(na2426_2), .IN1(na48_1), .IN2(1'b1), .IN3(~na33_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x77y84     80'h00_0078_00_0000_0C66_605C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2428_1 ( .OUT(na2428_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na36_1), .IN8(na35_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2428_4 ( .OUT(na2428_2), .IN1(1'b0), .IN2(na2413_2), .IN3(~na2409_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x82y97     80'h00_0018_00_0000_0EEE_0ADE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2429_1 ( .OUT(na2429_1), .IN1(na2430_1), .IN2(na2431_1), .IN3(~na57_2), .IN4(na61_1), .IN5(na2430_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x83y97     80'h00_0078_00_0000_0C88_5A8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2430_1 ( .OUT(na2430_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na11_1), .IN6(1'b1), .IN7(~na66_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2430_4 ( .OUT(na2430_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1001_1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y96     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2431_1 ( .OUT(na2431_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2220_2), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y95     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2432_1 ( .OUT(na2432_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1009_2), .IN6(~na2962_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y98     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2436_4 ( .OUT(na2436_2), .IN1(1'b1), .IN2(~na1084_1), .IN3(1'b1), .IN4(~na1083_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y68     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2438_1 ( .OUT(na2438_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3175_2), .IN7(1'b0), .IN8(na45_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x83y102     80'h00_0018_00_0000_0EEE_A5EE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2439_1 ( .OUT(na2439_1), .IN1(na2441_1), .IN2(na83_1), .IN3(na2440_1), .IN4(na2444_2), .IN5(~na2443_2), .IN6(1'b0), .IN7(na2440_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x82y99     80'h00_0078_00_0000_0C88_4FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2440_1 ( .OUT(na2440_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na66_2), .IN8(na69_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2440_4 ( .OUT(na2440_2), .IN1(na2221_1), .IN2(1'b1), .IN3(1'b1), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y99     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2441_1 ( .OUT(na2441_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(1'b1), .IN8(na69_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x83y99     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2443_4 ( .OUT(na2443_2), .IN1(~na1011_2), .IN2(1'b0), .IN3(~na2987_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y104     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2444_4 ( .OUT(na2444_2), .IN1(1'b1), .IN2(na1002_1), .IN3(1'b1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x82y86     80'h00_0018_00_0000_0EEE_E0CD
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2445_1 ( .OUT(na2445_1), .IN1(~na91_2), .IN2(na93_1), .IN3(1'b0), .IN4(na2447_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3177_2),
                      .IN8(na2446_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x88y92     80'h00_0078_00_0000_0C88_5CCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2446_1 ( .OUT(na2446_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(~na66_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2446_4 ( .OUT(na2446_2), .IN1(1'b1), .IN2(na1003_1), .IN3(1'b1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y90     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2447_1 ( .OUT(na2447_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2222_2), .IN6(1'b1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y89     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2448_1 ( .OUT(na2448_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1012_2), .IN6(~na85_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x82y88     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2450_4 ( .OUT(na2450_2), .IN1(na48_2), .IN2(na23_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y88     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2451_1 ( .OUT(na2451_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na48_1), .IN6(na23_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x84y84     80'h00_0018_00_0000_0EEE_30EE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2453_1 ( .OUT(na2453_1), .IN1(na103_1), .IN2(na2454_2), .IN3(na2457_1), .IN4(na2455_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(~na2456_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y86     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2454_4 ( .OUT(na2454_2), .IN1(na94_2), .IN2(na2989_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y88     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2455_1 ( .OUT(na2455_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2223_1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x86y86     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2456_4 ( .OUT(na2456_2), .IN1(~na82_1), .IN2(~na1013_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y91     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2457_1 ( .OUT(na2457_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1004_1), .IN7(1'b1), .IN8(na65_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x85y78     80'h00_0018_00_0000_0EEE_0CDE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2458_1 ( .OUT(na2458_1), .IN1(na2460_2), .IN2(na2459_1), .IN3(~na109_2), .IN4(na111_1), .IN5(1'b0), .IN6(na2459_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x87y86     80'h00_0078_00_0000_0C88_5C8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2459_1 ( .OUT(na2459_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na105_1), .IN7(~na66_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2459_4 ( .OUT(na2459_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1005_1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y81     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2460_4 ( .OUT(na2460_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2224_2), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y80     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2461_1 ( .OUT(na2461_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1014_2), .IN6(~na105_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x90y70     80'h00_0018_00_0000_0EEE_0CDE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2463_1 ( .OUT(na2463_1), .IN1(na119_1), .IN2(na2464_1), .IN3(~na120_2), .IN4(na2465_1), .IN5(1'b0), .IN6(na2464_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y80     80'h00_0078_00_0000_0C88_5ACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2464_1 ( .OUT(na2464_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na112_1), .IN6(1'b1), .IN7(~na66_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2464_4 ( .OUT(na2464_2), .IN1(na1006_1), .IN2(1'b1), .IN3(1'b1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y74     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2465_1 ( .OUT(na2465_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2225_1), .IN6(1'b1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y75     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2467_1 ( .OUT(na2467_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1015_2), .IN8(~na2996_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x88y82     80'h00_0018_00_0000_0888_7B75
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2469_1 ( .OUT(na2469_1), .IN1(~na127_1), .IN2(1'b0), .IN3(~na2226_2), .IN4(~na65_1), .IN5(na2472_1), .IN6(~na104_2), .IN7(~na1007_1),
                      .IN8(~na65_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y79     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2472_1 ( .OUT(na2472_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1016_2), .IN8(~na2997_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x85y77     80'h00_0018_00_0000_0EEE_DCEA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2473_1 ( .OUT(na2473_1), .IN1(na133_1), .IN2(1'b0), .IN3(na2478_2), .IN4(na2475_2), .IN5(1'b0), .IN6(na3178_2), .IN7(~na2477_1),
                      .IN8(na2474_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y82     80'h00_0078_00_0000_0C88_5ACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2474_1 ( .OUT(na2474_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na128_1), .IN6(1'b1), .IN7(~na66_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2474_4 ( .OUT(na2474_2), .IN1(1'b1), .IN2(na2227_1), .IN3(1'b1), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y80     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2475_4 ( .OUT(na2475_2), .IN1(na128_2), .IN2(1'b1), .IN3(na2988_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x88y79     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2477_1 ( .OUT(na2477_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1017_2), .IN6(1'b0), .IN7(~na2987_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y85     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2478_4 ( .OUT(na2478_2), .IN1(1'b1), .IN2(na2984_2), .IN3(1'b1), .IN4(na1008_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y84     80'h00_0018_00_0000_0EEE_C0ED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2479_1 ( .OUT(na2479_1), .IN1(~na139_1), .IN2(na2480_1), .IN3(na2481_2), .IN4(na137_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y86     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2480_1 ( .OUT(na2480_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1664_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y81     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2481_4 ( .OUT(na2481_2), .IN1(na82_1), .IN2(1'b1), .IN3(na929_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y94     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2482_1 ( .OUT(na2482_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1625_1), .IN6(1'b1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x97y92     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2484_4 ( .OUT(na2484_2), .IN1(~na82_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na1665_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x96y91     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2485_1 ( .OUT(na2485_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na747_1), .IN6(1'b1), .IN7(1'b1), .IN8(na65_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2485_4 ( .OUT(na2485_2), .IN1(na82_1), .IN2(1'b1), .IN3(1'b1), .IN4(na930_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y85     80'h00_0018_00_0000_0EEE_A0EB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2486_1 ( .OUT(na2486_1), .IN1(na149_1), .IN2(~na151_1), .IN3(na150_1), .IN4(na148_1), .IN5(1'b0), .IN6(1'b0), .IN7(na150_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x96y77     80'h00_0018_00_0000_0EEE_ACCD
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2489_1 ( .OUT(na2489_1), .IN1(~na156_1), .IN2(na155_1), .IN3(1'b0), .IN4(na2491_1), .IN5(1'b0), .IN6(na153_2), .IN7(na157_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y82     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2491_1 ( .OUT(na2491_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na932_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y77     80'h00_0018_00_0000_0888_F121
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2492_1 ( .OUT(na2492_1), .IN1(~na2493_2), .IN2(~na2495_1), .IN3(na2494_1), .IN4(~na163_1), .IN5(~na162_1), .IN6(~na2495_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y87     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2493_4 ( .OUT(na2493_2), .IN1(1'b1), .IN2(1'b1), .IN3(na763_1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x98y79     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2494_1 ( .OUT(na2494_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na82_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na1668_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x95y80     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2495_1 ( .OUT(na2495_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1628_2), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2495_4 ( .OUT(na2495_2), .IN1(na82_1), .IN2(1'b1), .IN3(1'b1), .IN4(na933_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y68     80'h00_0018_00_0000_0888_1325
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2497_1 ( .OUT(na2497_1), .IN1(~na169_1), .IN2(1'b1), .IN3(na2499_1), .IN4(~na2500_1), .IN5(1'b1), .IN6(~na168_1), .IN7(~na2498_2),
                      .IN8(~na2500_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y79     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2498_4 ( .OUT(na2498_2), .IN1(1'b1), .IN2(na2984_2), .IN3(1'b1), .IN4(na768_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x98y71     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2499_1 ( .OUT(na2499_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na82_2), .IN6(~na1669_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y74     80'h00_0078_00_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2500_1 ( .OUT(na2500_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1629_1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2500_4 ( .OUT(na2500_2), .IN1(na934_1), .IN2(1'b1), .IN3(na2987_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y71     80'h00_0018_00_0000_0EEE_CAEE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2502_1 ( .OUT(na2502_1), .IN1(na2504_1), .IN2(na173_1), .IN3(na175_1), .IN4(na2503_1), .IN5(na2504_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na2503_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x96y76     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2503_1 ( .OUT(na2503_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1630_2), .IN6(1'b1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2503_4 ( .OUT(na2503_2), .IN1(na82_2), .IN2(na1670_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y75     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2504_1 ( .OUT(na2504_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na770_1), .IN8(na65_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2504_4 ( .OUT(na2504_2), .IN1(na82_1), .IN2(1'b1), .IN3(1'b1), .IN4(na935_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y76     80'h00_0018_00_0000_0EEE_0EDE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2507_1 ( .OUT(na2507_1), .IN1(na181_1), .IN2(na178_1), .IN3(~na2509_2), .IN4(na2510_1), .IN5(na180_1), .IN6(na178_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x98y75     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2509_4 ( .OUT(na2509_2), .IN1(~na82_2), .IN2(1'b0), .IN3(~na1671_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y78     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2510_1 ( .OUT(na2510_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na773_1), .IN8(na65_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x84y104     80'h00_0018_00_0000_0888_3321
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2512_1 ( .OUT(na2512_1), .IN1(~na189_1), .IN2(~na2515_1), .IN3(na2514_1), .IN4(~na2513_2), .IN5(1'b1), .IN6(~na2515_2), .IN7(1'b1),
                      .IN8(~na188_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y100     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2513_4 ( .OUT(na2513_2), .IN1(1'b1), .IN2(na832_1), .IN3(1'b1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x90y103     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2514_1 ( .OUT(na2514_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na829_2), .IN6(1'b0), .IN7(~na2988_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y100     80'h00_0078_00_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2515_1 ( .OUT(na2515_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1658_2), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2515_4 ( .OUT(na2515_2), .IN1(na939_1), .IN2(1'b1), .IN3(na2987_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x85y97     80'h00_0018_00_0000_0EEE_EACE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2517_1 ( .OUT(na2517_1), .IN1(na194_1), .IN2(na195_2), .IN3(1'b0), .IN4(na2519_2), .IN5(na193_1), .IN6(1'b0), .IN7(na3179_2),
                      .IN8(na2518_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y98     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2518_1 ( .OUT(na2518_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(na833_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2518_4 ( .OUT(na2518_2), .IN1(na82_1), .IN2(1'b1), .IN3(1'b1), .IN4(na940_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y94     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2519_4 ( .OUT(na2519_2), .IN1(1'b1), .IN2(na1659_1), .IN3(1'b1), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x92y96     80'h00_0018_00_0000_0EEE_E03E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2521_1 ( .OUT(na2521_1), .IN1(na199_1), .IN2(na2523_2), .IN3(1'b0), .IN4(~na201_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2522_1),
                      .IN8(na200_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y99     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2522_1 ( .OUT(na2522_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na839_2), .IN6(1'b1), .IN7(na2988_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y96     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2523_4 ( .OUT(na2523_2), .IN1(na82_1), .IN2(na941_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x100y85     80'h00_0018_00_0000_0EEE_CEAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2524_1 ( .OUT(na2524_1), .IN1(na2525_1), .IN2(na2526_2), .IN3(na205_1), .IN4(1'b0), .IN5(na2525_2), .IN6(na2526_1), .IN7(1'b0),
                      .IN8(na207_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x101y91     80'h00_0078_00_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2525_1 ( .OUT(na2525_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na842_2), .IN6(1'b1), .IN7(na2988_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2525_4 ( .OUT(na2525_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1661_1), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x99y88     80'h00_0078_00_0000_0C88_CA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2526_1 ( .OUT(na2526_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(1'b1), .IN8(na942_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2526_4 ( .OUT(na2526_2), .IN1(1'b1), .IN2(1'b1), .IN3(na844_1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y88     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2529_1 ( .OUT(na2529_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na845_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2529_4 ( .OUT(na2529_2), .IN1(na943_1), .IN2(1'b1), .IN3(na2987_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y97     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2531_1 ( .OUT(na2531_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1663_1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x107y101     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2533_4 ( .OUT(na2533_2), .IN1(~na847_2), .IN2(~na2989_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x100y96     80'h00_0078_00_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2534_1 ( .OUT(na2534_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na848_1), .IN7(1'b1), .IN8(na65_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2534_4 ( .OUT(na2534_2), .IN1(na82_1), .IN2(na944_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x88y96     80'h00_0018_00_0000_0EEE_D0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2535_1 ( .OUT(na2535_1), .IN1(1'b0), .IN2(na223_1), .IN3(na2537_1), .IN4(na2536_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na225_1),
                      .IN8(na224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y94     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2536_1 ( .OUT(na2536_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(na2228_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y93     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2537_1 ( .OUT(na2537_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na945_1), .IN6(1'b1), .IN7(na2987_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x89y105     80'h00_0018_00_0000_0EEE_AACD
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2538_1 ( .OUT(na2538_1), .IN1(~na230_1), .IN2(na229_1), .IN3(1'b0), .IN4(na2540_2), .IN5(na231_1), .IN6(1'b0), .IN7(na227_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y104     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2540_4 ( .OUT(na2540_2), .IN1(na82_1), .IN2(na946_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y98     80'h00_0018_00_0000_0EEE_CAEE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2541_1 ( .OUT(na2541_1), .IN1(na2543_1), .IN2(na235_1), .IN3(na237_1), .IN4(na2542_1), .IN5(na2543_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na2542_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y98     80'h00_0078_00_0000_0C88_F8CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2542_1 ( .OUT(na2542_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(na2230_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2542_4 ( .OUT(na2542_2), .IN1(1'b1), .IN2(na908_2), .IN3(1'b1), .IN4(na65_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x91y95     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2543_1 ( .OUT(na2543_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na947_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2543_4 ( .OUT(na2543_2), .IN1(na911_1), .IN2(1'b1), .IN3(1'b1), .IN4(na65_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y90     80'h00_0018_00_0000_0888_1325
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2546_1 ( .OUT(na2546_1), .IN1(~na3181_2), .IN2(1'b1), .IN3(na2548_2), .IN4(~na2547_1), .IN5(1'b1), .IN6(~na243_1), .IN7(~na242_1),
                      .IN8(~na2549_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y88     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2547_1 ( .OUT(na2547_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2984_2), .IN7(1'b1), .IN8(na917_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x92y89     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2548_4 ( .OUT(na2548_2), .IN1(~na2231_1), .IN2(1'b0), .IN3(~na2988_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y90     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2549_1 ( .OUT(na2549_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na912_2), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2549_4 ( .OUT(na2549_2), .IN1(na82_1), .IN2(na948_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x91y85     80'h00_0018_00_0000_0EEE_A0ED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2551_1 ( .OUT(na2551_1), .IN1(~na248_1), .IN2(na247_1), .IN3(na245_1), .IN4(na2553_1), .IN5(1'b0), .IN6(1'b0), .IN7(na249_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y86     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2553_1 ( .OUT(na2553_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na949_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x94y78     80'h00_0018_00_0000_0EEE_AEAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2554_1 ( .OUT(na2554_1), .IN1(na253_1), .IN2(na2555_1), .IN3(na2556_1), .IN4(1'b0), .IN5(na255_1), .IN6(na2555_2), .IN7(na2556_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y84     80'h00_0078_00_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2555_1 ( .OUT(na2555_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na921_2), .IN6(1'b1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2555_4 ( .OUT(na2555_2), .IN1(na82_2), .IN2(na2233_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x96y83     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2556_1 ( .OUT(na2556_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2983_2), .IN8(na924_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2556_4 ( .OUT(na2556_2), .IN1(na82_1), .IN2(na950_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x93y73     80'h00_0018_00_0000_0EEE_0EBE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2559_1 ( .OUT(na2559_1), .IN1(na2562_1), .IN2(na258_1), .IN3(na261_1), .IN4(~na2561_2), .IN5(na260_1), .IN6(na258_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x94y86     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2561_4 ( .OUT(na2561_2), .IN1(~na82_2), .IN2(1'b0), .IN3(~na2234_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y79     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2562_1 ( .OUT(na2562_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na926_1), .IN7(1'b1), .IN8(na65_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x94y80     80'h00_0018_00_0000_0EEE_EAEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2564_1 ( .OUT(na2564_1), .IN1(1'b0), .IN2(na265_1), .IN3(na267_1), .IN4(na2566_1), .IN5(na3182_2), .IN6(1'b0), .IN7(na2565_2),
                      .IN8(na2566_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x96y81     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2565_1 ( .OUT(na2565_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na927_2), .IN6(1'b1), .IN7(1'b1), .IN8(na65_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2565_4 ( .OUT(na2565_2), .IN1(na82_2), .IN2(1'b1), .IN3(na2235_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x94y84     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2566_1 ( .OUT(na2566_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2983_2), .IN8(na928_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2566_4 ( .OUT(na2566_2), .IN1(na82_1), .IN2(na952_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y101     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2570_1 ( .OUT(na2570_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na589_1), .IN6(na493_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y101     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2571_1 ( .OUT(na2571_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3049_2), .IN8(~na653_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x86y102     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2572_1 ( .OUT(na2572_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na654_1), .IN6(1'b1), .IN7(na2987_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2572_4 ( .OUT(na2572_2), .IN1(na82_2), .IN2(na558_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x86y100     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2573_1 ( .OUT(na2573_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na430_2), .IN6(na470_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y92     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2575_1 ( .OUT(na2575_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na655_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2575_4 ( .OUT(na2575_2), .IN1(na82_2), .IN2(1'b1), .IN3(na559_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y90     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2576_1 ( .OUT(na2576_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3156_2), .IN5(1'b0), .IN6(na495_1), .IN7(1'b0), .IN8(na591_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y83     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2578_1 ( .OUT(na2578_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na656_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2578_4 ( .OUT(na2578_2), .IN1(na82_2), .IN2(1'b1), .IN3(na560_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y79     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2579_1 ( .OUT(na2579_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na592_1), .IN6(na496_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y74     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2581_1 ( .OUT(na2581_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na657_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2581_4 ( .OUT(na2581_2), .IN1(na82_2), .IN2(na561_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y74     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2582_1 ( .OUT(na2582_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na497_2), .IN6(na593_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y70     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2584_1 ( .OUT(na2584_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(1'b1), .IN8(na658_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2584_4 ( .OUT(na2584_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na562_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x98y67     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2585_1 ( .OUT(na2585_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na498_2), .IN6(na594_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x94y70     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2587_1 ( .OUT(na2587_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na659_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2587_4 ( .OUT(na2587_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na563_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y70     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2588_1 ( .OUT(na2588_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na595_2), .IN8(na499_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x95y72     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2590_1 ( .OUT(na2590_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na660_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2590_4 ( .OUT(na2590_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na564_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y72     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2591_1 ( .OUT(na2591_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3156_2), .IN5(na500_1), .IN6(1'b0), .IN7(na596_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x107y91     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2593_1 ( .OUT(na2593_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(1'b1), .IN8(na565_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2593_4 ( .OUT(na2593_2), .IN1(na82_1), .IN2(1'b1), .IN3(1'b1), .IN4(na661_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y91     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2594_1 ( .OUT(na2594_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na3156_2), .IN5(na597_2), .IN6(1'b0), .IN7(na501_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x102y100     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2596_1 ( .OUT(na2596_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na662_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2596_4 ( .OUT(na2596_2), .IN1(na82_2), .IN2(na566_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y100     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2597_1 ( .OUT(na2597_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na438_2), .IN8(na478_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x110y88     80'h00_0078_00_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2599_1 ( .OUT(na2599_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(1'b1), .IN8(na567_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2599_4 ( .OUT(na2599_2), .IN1(na82_1), .IN2(1'b1), .IN3(1'b1), .IN4(na663_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y83     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2600_1 ( .OUT(na2600_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na599_1), .IN8(na503_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y80     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2602_1 ( .OUT(na2602_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na664_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2602_4 ( .OUT(na2602_2), .IN1(na82_2), .IN2(na568_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y79     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2603_1 ( .OUT(na2603_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3156_2), .IN5(na504_2), .IN6(1'b0), .IN7(na600_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y77     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2605_1 ( .OUT(na2605_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na665_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2605_4 ( .OUT(na2605_2), .IN1(na82_2), .IN2(1'b1), .IN3(na569_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x112y80     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2606_1 ( .OUT(na2606_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na601_1), .IN8(na505_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x106y71     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2608_1 ( .OUT(na2608_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na570_1), .IN6(1'b1), .IN7(na2988_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2608_4 ( .OUT(na2608_2), .IN1(na666_1), .IN2(1'b1), .IN3(na2987_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y69     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2609_1 ( .OUT(na2609_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na602_2), .IN6(na506_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y75     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2611_1 ( .OUT(na2611_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(1'b1), .IN7(1'b1), .IN8(na571_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2611_4 ( .OUT(na2611_2), .IN1(na82_1), .IN2(1'b1), .IN3(na667_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y72     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2612_1 ( .OUT(na2612_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3156_2), .IN5(1'b0), .IN6(na507_1), .IN7(1'b0), .IN8(na603_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x106y76     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2614_1 ( .OUT(na2614_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na668_1), .IN6(1'b1), .IN7(na2987_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2614_4 ( .OUT(na2614_2), .IN1(na82_2), .IN2(na572_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y72     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2615_1 ( .OUT(na2615_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na604_2), .IN8(na508_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x109y86     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2617_1 ( .OUT(na2617_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(na573_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2617_4 ( .OUT(na2617_2), .IN1(na669_2), .IN2(1'b1), .IN3(na2987_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y85     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2618_1 ( .OUT(na2618_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na509_1), .IN6(na605_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x106y80     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2620_1 ( .OUT(na2620_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na670_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2620_4 ( .OUT(na2620_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na574_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y81     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2621_1 ( .OUT(na2621_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3156_2), .IN5(1'b0), .IN6(na510_2), .IN7(1'b0), .IN8(na606_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y103     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2623_1 ( .OUT(na2623_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na671_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2623_4 ( .OUT(na2623_2), .IN1(na82_2), .IN2(1'b1), .IN3(na575_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y106     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2624_1 ( .OUT(na2624_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3156_2), .IN5(1'b0), .IN6(na607_1), .IN7(1'b0), .IN8(na511_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y94     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2626_1 ( .OUT(na2626_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na672_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2626_4 ( .OUT(na2626_2), .IN1(na82_2), .IN2(1'b1), .IN3(na576_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x111y93     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2627_1 ( .OUT(na2627_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na3156_2), .IN5(na608_2), .IN6(1'b0), .IN7(na512_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x100y99     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2629_1 ( .OUT(na2629_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(na577_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2629_4 ( .OUT(na2629_2), .IN1(na673_2), .IN2(1'b1), .IN3(na2987_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x104y101     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2630_1 ( .OUT(na2630_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na3156_2), .IN5(na3052_2), .IN6(1'b0), .IN7(na513_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x112y88     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2632_1 ( .OUT(na2632_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na674_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2632_4 ( .OUT(na2632_2), .IN1(na82_2), .IN2(na578_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x115y89     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2633_1 ( .OUT(na2633_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3156_2), .IN5(na3023_2), .IN6(1'b0), .IN7(na490_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x110y75     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2635_1 ( .OUT(na2635_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na675_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2635_4 ( .OUT(na2635_2), .IN1(na82_2), .IN2(na579_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x109y78     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2636_1 ( .OUT(na2636_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3156_2), .IN5(1'b0), .IN6(na515_2), .IN7(1'b0), .IN8(na611_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y99     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2638_1 ( .OUT(na2638_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na676_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2638_4 ( .OUT(na2638_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na580_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x103y97     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2639_1 ( .OUT(na2639_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na452_2), .IN8(na492_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y92     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2641_1 ( .OUT(na2641_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(na581_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2641_4 ( .OUT(na2641_2), .IN1(na82_1), .IN2(na677_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y93     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2642_1 ( .OUT(na2642_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na517_1), .IN8(na461_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y104     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2644_1 ( .OUT(na2644_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na678_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2644_4 ( .OUT(na2644_2), .IN1(na82_2), .IN2(na582_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y102     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2645_1 ( .OUT(na2645_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na518_1), .IN6(na462_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y100     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2647_1 ( .OUT(na2647_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na679_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2647_4 ( .OUT(na2647_2), .IN1(na82_2), .IN2(na583_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y100     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2648_1 ( .OUT(na2648_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na615_1), .IN8(na519_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y91     80'h00_0078_00_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2650_1 ( .OUT(na2650_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(na680_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2650_4 ( .OUT(na2650_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na584_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y89     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2651_1 ( .OUT(na2651_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3156_2), .IN5(1'b0), .IN6(na616_2), .IN7(1'b0), .IN8(na520_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y85     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2653_1 ( .OUT(na2653_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(na585_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2653_4 ( .OUT(na2653_2), .IN1(na82_1), .IN2(1'b1), .IN3(na681_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x108y86     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2654_1 ( .OUT(na2654_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na521_2), .IN6(na617_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x106y73     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2656_1 ( .OUT(na2656_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na682_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2656_4 ( .OUT(na2656_2), .IN1(na82_2), .IN2(1'b1), .IN3(na586_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x110y74     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2657_1 ( .OUT(na2657_1), .IN1(~na1087_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na618_2), .IN8(na522_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x99y72     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2659_1 ( .OUT(na2659_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_2), .IN6(na587_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2659_4 ( .OUT(na2659_2), .IN1(na82_1), .IN2(1'b1), .IN3(na683_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y72     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2660_1 ( .OUT(na2660_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3156_2), .IN5(1'b0), .IN6(na467_2), .IN7(1'b0), .IN8(na523_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x102y75     80'h00_0078_00_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2662_1 ( .OUT(na2662_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(na684_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2662_4 ( .OUT(na2662_2), .IN1(na82_2), .IN2(1'b1), .IN3(1'b1), .IN4(na588_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y78     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2663_1 ( .OUT(na2663_1), .IN1(na1087_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3043_2), .IN6(na468_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y73     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2668_4 ( .OUT(na2668_2), .IN1(1'b0), .IN2(na713_1), .IN3(1'b0), .IN4(na697_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x122y85     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2669_1 ( .OUT(na2669_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na702_1), .IN5(1'b0), .IN6(~na3136_2), .IN7(1'b0), .IN8(~na1039_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y85     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2670_4 ( .OUT(na2670_2), .IN1(na1045_1), .IN2(na704_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x124y79     80'h00_0078_00_0000_0C88_C3A5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2671_1 ( .OUT(na2671_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na704_2), .IN7(1'b1), .IN8(na702_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2671_4 ( .OUT(na2671_2), .IN1(~na703_2), .IN2(1'b1), .IN3(na706_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x124y85     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2672_1 ( .OUT(na2672_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1035_1), .IN8(na702_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y86     80'h00_0060_00_0000_0C06_FFC3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2677_4 ( .OUT(na2677_2), .IN1(1'b0), .IN2(~na704_2), .IN3(1'b0), .IN4(na1039_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y68     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2678_4 ( .OUT(na2678_2), .IN1(na1458_1), .IN2(1'b0), .IN3(1'b0), .IN4(na697_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y73     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2680_1 ( .OUT(na2680_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na709_1), .IN8(na697_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y74     80'h00_0060_00_0000_0C06_FFA3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2682_4 ( .OUT(na2682_2), .IN1(1'b0), .IN2(~na713_1), .IN3(na709_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y70     80'h00_0018_00_0000_0C66_5A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2684_1 ( .OUT(na2684_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na725_2), .IN6(1'b0), .IN7(~na724_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y65     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2685_1 ( .OUT(na2685_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na724_1), .IN8(~na2693_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y69     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2686_4 ( .OUT(na2686_2), .IN1(~na725_2), .IN2(1'b0), .IN3(1'b0), .IN4(na729_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y80     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2688_1 ( .OUT(na2688_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3069_2), .IN8(na702_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y75     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2690_4 ( .OUT(na2690_2), .IN1(~na737_1), .IN2(1'b0), .IN3(1'b0), .IN4(na729_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x109y85     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2691_1 ( .OUT(na2691_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2371_1), .IN7(1'b0), .IN8(na308_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x124y70     80'h00_0078_00_0000_0C66_90C9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2693_1 ( .OUT(na2693_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na717_1), .IN8(~na729_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2693_4 ( .OUT(na2693_2), .IN1(na3064_2), .IN2(~na704_2), .IN3(1'b0), .IN4(na729_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x122y67     80'h00_0078_00_0000_0C88_AAC3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2694_1 ( .OUT(na2694_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na725_2), .IN6(1'b1), .IN7(na717_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2694_4 ( .OUT(na2694_2), .IN1(1'b1), .IN2(~na720_1), .IN3(1'b1), .IN4(na729_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y63     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2696_4 ( .OUT(na2696_2), .IN1(1'b0), .IN2(na722_1), .IN3(na724_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x104y91     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2697_1 ( .OUT(na2697_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na313_1), .IN6(1'b0), .IN7(1'b0), .IN8(na2372_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x106y81     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2698_4 ( .OUT(na2698_2), .IN1(na2373_1), .IN2(1'b0), .IN3(1'b0), .IN4(na318_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x119y72     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2699_1 ( .OUT(na2699_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na703_2), .IN6(1'b0), .IN7(1'b0), .IN8(na729_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y76     80'h00_0060_00_0000_0C06_FF3A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2700_4 ( .OUT(na2700_2), .IN1(na737_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na702_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x104y77     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2701_1 ( .OUT(na2701_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2374_1), .IN7(na323_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x105y79     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2702_4 ( .OUT(na2702_2), .IN1(na328_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2375_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x107y67     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2703_1 ( .OUT(na2703_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2376_1), .IN7(na333_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x104y75     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2704_4 ( .OUT(na2704_2), .IN1(1'b0), .IN2(na338_1), .IN3(na2377_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x101y73     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2705_1 ( .OUT(na2705_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2378_1), .IN6(1'b0), .IN7(1'b0), .IN8(na343_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x126y108     80'h00_0078_00_0000_0C66_ACA9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2706_1 ( .OUT(na2706_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2724_2), .IN7(na797_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2706_4 ( .OUT(na2706_2), .IN1(~na800_1), .IN2(na779_1), .IN3(na780_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y97     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2707_4 ( .OUT(na2707_2), .IN1(1'b0), .IN2(na3197_2), .IN3(na791_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x120y101     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2712_4 ( .OUT(na2712_2), .IN1(1'b0), .IN2(na779_1), .IN3(na780_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x123y94     80'h00_0078_00_0000_0C88_C32F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2714_1 ( .OUT(na2714_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na779_1), .IN7(1'b1), .IN8(na781_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2714_4 ( .OUT(na2714_2), .IN1(1'b1), .IN2(1'b1), .IN3(na783_2), .IN4(~na2722_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x121y90     80'h00_0078_00_0000_0C66_90A9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2716_1 ( .OUT(na2716_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na780_2), .IN8(~na1051_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2716_4 ( .OUT(na2716_2), .IN1(na1059_1), .IN2(~na1063_1), .IN3(na1061_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x125y101     80'h00_0078_00_0000_0C66_60A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2718_1 ( .OUT(na2718_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na791_1), .IN8(na1461_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2718_4 ( .OUT(na2718_2), .IN1(na795_2), .IN2(na796_1), .IN3(na1462_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y106     80'h00_0060_00_0000_0C06_FF3A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2719_4 ( .OUT(na2719_2), .IN1(na804_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na806_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x126y96     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2720_1 ( .OUT(na2720_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na786_1), .IN6(na3197_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x124y99     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2721_4 ( .OUT(na2721_2), .IN1(1'b0), .IN2(na3197_2), .IN3(1'b0), .IN4(~na1461_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x124y90     80'h00_0078_00_0000_0C66_AC90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2722_1 ( .OUT(na2722_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2716_2), .IN7(na3102_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2722_4 ( .OUT(na2722_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1061_1), .IN4(na1065_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y100     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2723_1 ( .OUT(na2723_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na797_1), .IN8(~na781_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x121y106     80'h00_0078_00_0000_0C66_A5C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2724_1 ( .OUT(na2724_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na778_1), .IN6(1'b0), .IN7(na797_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2724_4 ( .OUT(na2724_2), .IN1(1'b0), .IN2(~na779_1), .IN3(1'b0), .IN4(na781_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x123y95     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2725_4 ( .OUT(na2725_2), .IN1(na800_1), .IN2(1'b0), .IN3(~na812_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x122y95     80'h00_0078_00_0000_0C66_3C90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2729_1 ( .OUT(na2729_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na802_1), .IN7(1'b0), .IN8(~na1051_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2729_4 ( .OUT(na2729_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na780_2), .IN4(na2722_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x122y106     80'h00_0018_00_0000_0C66_C300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2730_1 ( .OUT(na2730_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na2724_2), .IN7(1'b0), .IN8(na806_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x110y94     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2731_4 ( .OUT(na2731_2), .IN1(1'b0), .IN2(1'b0), .IN3(na348_1), .IN4(na2379_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y101     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2733_1 ( .OUT(na2733_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2724_2), .IN7(na2729_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y107     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2734_4 ( .OUT(na2734_2), .IN1(na804_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2706_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x108y92     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2736_1 ( .OUT(na2736_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2380_1), .IN6(1'b0), .IN7(na353_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x96y103     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2737_4 ( .OUT(na2737_2), .IN1(na2381_1), .IN2(1'b0), .IN3(na358_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y98     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2738_1 ( .OUT(na2738_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na800_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na781_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x119y90     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2739_4 ( .OUT(na2739_2), .IN1(1'b0), .IN2(1'b0), .IN3(na812_1), .IN4(na781_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x100y98     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2740_1 ( .OUT(na2740_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2382_1), .IN6(1'b0), .IN7(1'b0), .IN8(na363_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x106y101     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2741_4 ( .OUT(na2741_2), .IN1(1'b0), .IN2(1'b0), .IN3(na368_1), .IN4(na2383_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y89     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2742_1 ( .OUT(na2742_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2384_1), .IN6(na373_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x109y85     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2743_4 ( .OUT(na2743_2), .IN1(1'b0), .IN2(na378_1), .IN3(na2385_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x106y101     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2744_1 ( .OUT(na2744_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2386_1), .IN7(1'b0), .IN8(na383_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x125y107     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2745_4 ( .OUT(na2745_2), .IN1(1'b0), .IN2(na879_2), .IN3(na878_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x125y109     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2746_1 ( .OUT(na2746_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2758_2), .IN8(~na868_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x116y107     80'h00_0078_00_0000_0C88_F835
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2748_1 ( .OUT(na2748_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2750_2), .IN6(na860_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2748_4 ( .OUT(na2748_2), .IN1(~na856_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na858_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x115y103     80'h00_0078_00_0000_0C66_A699
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2750_1 ( .OUT(na2750_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na856_1), .IN6(na1067_1), .IN7(na2757_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2750_4 ( .OUT(na2750_2), .IN1(na1071_1), .IN2(~na3149_2), .IN3(~na1069_1), .IN4(na1075_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x114y103     80'h00_0078_00_0000_0C66_CA90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2751_1 ( .OUT(na2751_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na856_1), .IN6(1'b0), .IN7(1'b0), .IN8(na858_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2751_4 ( .OUT(na2751_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1069_1), .IN4(na1081_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x117y105     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2756_4 ( .OUT(na2756_2), .IN1(~na856_1), .IN2(na1067_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x116y105     80'h00_0078_00_0000_0C66_09C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2757_1 ( .OUT(na2757_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na870_2), .IN6(na1077_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2757_4 ( .OUT(na2757_2), .IN1(~na1071_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1075_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x118y111     80'h00_0078_00_0000_0C66_CAA6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2758_1 ( .OUT(na2758_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1465_1), .IN6(1'b0), .IN7(1'b0), .IN8(na868_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2758_4 ( .OUT(na2758_2), .IN1(na875_1), .IN2(na876_1), .IN3(na874_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x121y107     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2759_1 ( .OUT(na2759_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3121_2), .IN6(1'b0), .IN7(na884_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x122y110     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2760_4 ( .OUT(na2760_2), .IN1(1'b0), .IN2(na863_1), .IN3(na2758_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x116y108     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2761_1 ( .OUT(na2761_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1465_1), .IN6(~na863_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x120y107     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2762_4 ( .OUT(na2762_2), .IN1(na856_1), .IN2(1'b0), .IN3(1'b0), .IN4(na882_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x113y107     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2763_1 ( .OUT(na2763_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na860_1), .IN7(1'b0), .IN8(na858_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x115y108     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2765_4 ( .OUT(na2765_2), .IN1(~na892_1), .IN2(1'b0), .IN3(1'b0), .IN4(na880_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x117y102     80'h00_0078_00_0000_0C88_CC33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2766_1 ( .OUT(na2766_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na860_1), .IN7(1'b1), .IN8(na882_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2766_4 ( .OUT(na2766_2), .IN1(1'b1), .IN2(~na883_1), .IN3(1'b1), .IN4(~na858_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x118y105     80'h00_0078_00_0000_0C66_C35C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2769_1 ( .OUT(na2769_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1067_1), .IN7(1'b0), .IN8(na882_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2769_4 ( .OUT(na2769_2), .IN1(1'b0), .IN2(na860_2), .IN3(~na2757_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x120y106     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2770_1 ( .OUT(na2770_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3121_2), .IN6(1'b0), .IN7(na878_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x96y97     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2771_4 ( .OUT(na2771_2), .IN1(1'b0), .IN2(na2387_1), .IN3(na388_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x118y106     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2773_1 ( .OUT(na2773_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na879_2), .IN7(na884_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x97y110     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2774_4 ( .OUT(na2774_2), .IN1(1'b0), .IN2(1'b0), .IN3(na393_1), .IN4(na2388_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x91y103     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2775_1 ( .OUT(na2775_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2389_1), .IN6(1'b0), .IN7(1'b0), .IN8(na398_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x120y105     80'h00_0060_00_0000_0C06_FF3A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2776_4 ( .OUT(na2776_2), .IN1(na892_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na858_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x114y106     80'h00_0018_00_0000_0C66_C300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2777_1 ( .OUT(na2777_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na860_1), .IN7(1'b0), .IN8(na880_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x93y93     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2778_4 ( .OUT(na2778_2), .IN1(1'b0), .IN2(na2390_1), .IN3(na403_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x99y91     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2779_1 ( .OUT(na2779_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2391_1), .IN6(1'b0), .IN7(na408_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x102y81     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2780_4 ( .OUT(na2780_2), .IN1(1'b0), .IN2(na413_1), .IN3(1'b0), .IN4(na2392_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x100y77     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2781_1 ( .OUT(na2781_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2393_1), .IN7(1'b0), .IN8(na418_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x102y85     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2782_4 ( .OUT(na2782_2), .IN1(na423_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2394_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x107y96     80'h00_0078_00_0000_0C66_6006
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2855_1 ( .OUT(na2855_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2363_1), .IN8(na268_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2855_4 ( .OUT(na2855_2), .IN1(na1085_1), .IN2(na2436_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y104     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2856_1 ( .OUT(na2856_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na273_1), .IN8(na2364_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x86y96     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2857_4 ( .OUT(na2857_2), .IN1(na2365_1), .IN2(1'b0), .IN3(na278_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y87     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2858_1 ( .OUT(na2858_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na283_1), .IN8(na2366_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x86y82     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2859_4 ( .OUT(na2859_2), .IN1(1'b0), .IN2(na2367_1), .IN3(1'b0), .IN4(na288_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x92y77     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2860_1 ( .OUT(na2860_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2368_1), .IN7(1'b0), .IN8(na293_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x90y81     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2861_4 ( .OUT(na2861_2), .IN1(na298_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2369_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x90y81     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2862_1 ( .OUT(na2862_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na303_1), .IN8(na2370_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x84y108     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2904_4 ( .OUT(na2904_2), .IN1(1'b1), .IN2(na2408_2), .IN3(na3152_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y110     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2905_1 ( .OUT(na2905_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1085_1), .IN6(na2408_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x84y102     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2906_1 ( .OUT(na2906_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1084_1), .IN7(na66_1), .IN8(na1083_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y110     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2908_4 ( .OUT(na2908_2), .IN1(na1085_1), .IN2(~na2408_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y89     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2909_1 ( .OUT(na2909_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3011_2), .IN8(na1010_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y86     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2912_1 ( .OUT(na2912_1), .IN1(1'b1), .IN2(~na3012_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1103_2), .IN8(na2986_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y102     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2918_4 ( .OUT(na2918_2), .IN1(1'b1), .IN2(~na1084_1), .IN3(1'b1), .IN4(na1010_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y84     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2922_1 ( .OUT(na2922_1), .IN1(1'b1), .IN2(na3012_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na66_1), .IN8(na2994_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x101y86     80'h00_0078_00_0000_0C88_4F13
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2923_1 ( .OUT(na2923_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na66_2), .IN8(na429_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2923_4 ( .OUT(na2923_2), .IN1(1'b1), .IN2(~na1090_2), .IN3(~na1089_2), .IN4(~na3157_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y81     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2925_1 ( .OUT(na2925_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2349_1), .IN7(~na2351_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x86y81     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2926_4 ( .OUT(na2926_2), .IN1(1'b1), .IN2(na2349_1), .IN3(na2351_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x84y78     80'h00_0018_00_0000_0EEE_3EED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2927_1 ( .OUT(na2927_1), .IN1(~na6_1), .IN2(na5_2), .IN3(na8_2), .IN4(na7_1), .IN5(na6_2), .IN6(na5_1), .IN7(1'b0), .IN8(~na7_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x81y89     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2930_1 ( .OUT(na2930_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1033_1), .IN6(na23_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x83y91     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2931_4 ( .OUT(na2931_2), .IN1(1'b0), .IN2(na1031_1), .IN3(na1018_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x79y110     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2933_1 ( .OUT(na2933_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na20_2), .IN6(1'b0), .IN7(1'b0), .IN8(na25_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x80y101     80'h00_0078_00_0000_0C88_F255
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2934_1 ( .OUT(na2934_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na20_1), .IN6(~na23_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2934_4 ( .OUT(na2934_2), .IN1(~na20_2), .IN2(1'b1), .IN3(~na2409_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x99y94     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2936_4 ( .OUT(na2936_2), .IN1(~na82_2), .IN2(~na774_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y94     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2937_1 ( .OUT(na2937_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(1'b1), .IN8(na937_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x102y95     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a2939_4 ( .OUT(na2939_2), .IN1(~na82_2), .IN2(~na820_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y92     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2940_1 ( .OUT(na2940_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na82_1), .IN6(1'b1), .IN7(1'b1), .IN8(na938_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y82     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2942_1 ( .OUT(na2942_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na702_1), .IN5(1'b0), .IN6(~na704_2), .IN7(1'b0), .IN8(~na700_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x118y107     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2950_4 ( .OUT(na2950_2), .IN1(1'b0), .IN2(na1067_1), .IN3(na2757_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x117y108     80'h00_0018_00_0000_0C66_5A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2951_1 ( .OUT(na2951_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na853_1), .IN6(1'b0), .IN7(~na877_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x107y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2952_4 ( .OUT(na2952_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1001_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2952_6 ( .RAM_O2(na2952_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2952_2), .COMP_OUT(1'b0) );
// C_///AND/      x111y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2953_4 ( .OUT(na2953_2), .IN1(1'b1), .IN2(na1002_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2953_6 ( .RAM_O2(na2953_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2953_2), .COMP_OUT(1'b0) );
// C_///AND/      x115y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2954_4 ( .OUT(na2954_2), .IN1(1'b1), .IN2(na1003_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2954_6 ( .RAM_O2(na2954_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2954_2), .COMP_OUT(1'b0) );
// C_///AND/      x119y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2955_4 ( .OUT(na2955_2), .IN1(1'b1), .IN2(na1004_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2955_6 ( .RAM_O2(na2955_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2955_2), .COMP_OUT(1'b0) );
// C_///AND/      x123y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2956_4 ( .OUT(na2956_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1005_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2956_6 ( .RAM_O2(na2956_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2956_2), .COMP_OUT(1'b0) );
// C_///AND/      x127y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2957_4 ( .OUT(na2957_2), .IN1(na1006_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2957_6 ( .RAM_O2(na2957_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2957_2), .COMP_OUT(1'b0) );
// C_///AND/      x131y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2958_4 ( .OUT(na2958_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1007_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2958_6 ( .RAM_O2(na2958_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2958_2), .COMP_OUT(1'b0) );
// C_///AND/      x135y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2959_4 ( .OUT(na2959_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1008_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a2959_6 ( .RAM_O2(na2959_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na2959_2), .COMP_OUT(1'b0) );
// C_////Bridge      x88y68     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2960_5 ( .OUT(na2960_2), .IN1(1'b0), .IN2(na2_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y84     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2961_5 ( .OUT(na2961_2), .IN1(1'b0), .IN2(na5_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y96     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2962_5 ( .OUT(na2962_2), .IN1(na11_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y91     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2963_5 ( .OUT(na2963_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na15_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2964_5 ( .OUT(na2964_2), .IN1(na18_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y106     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2965_5 ( .OUT(na2965_2), .IN1(na20_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y103     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2966_5 ( .OUT(na2966_2), .IN1(na20_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y78     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2967_5 ( .OUT(na2967_2), .IN1(1'b0), .IN2(na23_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y108     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2968_5 ( .OUT(na2968_2), .IN1(1'b0), .IN2(na23_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y95     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2969_5 ( .OUT(na2969_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na23_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y79     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2970_5 ( .OUT(na2970_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na27_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y93     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2971_5 ( .OUT(na2971_2), .IN1(1'b0), .IN2(1'b0), .IN3(na33_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y83     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2972_5 ( .OUT(na2972_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na35_1) );
// C_////Bridge      x84y92     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2973_5 ( .OUT(na2973_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na42_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2974_5 ( .OUT(na2974_2), .IN1(na42_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y65     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2975_5 ( .OUT(na2975_2), .IN1(na42_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2976_5 ( .OUT(na2976_2), .IN1(na42_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2977_5 ( .OUT(na2977_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na43_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y69     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2978_5 ( .OUT(na2978_2), .IN1(na48_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2979_5 ( .OUT(na2979_2), .IN1(na48_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y71     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2980_5 ( .OUT(na2980_2), .IN1(na48_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2981_5 ( .OUT(na2981_2), .IN1(1'b0), .IN2(na49_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y84     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2982_5 ( .OUT(na2982_2), .IN1(1'b0), .IN2(na62_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y83     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2983_5 ( .OUT(na2983_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na65_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y82     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2984_5 ( .OUT(na2984_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na65_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2985_5 ( .OUT(na2985_2), .IN1(1'b0), .IN2(1'b0), .IN3(na66_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y90     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2986_5 ( .OUT(na2986_2), .IN1(1'b0), .IN2(1'b0), .IN3(na66_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2987_5 ( .OUT(na2987_2), .IN1(na82_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2988_5 ( .OUT(na2988_2), .IN1(na82_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y94     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2989_5 ( .OUT(na2989_2), .IN1(na82_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2990_5 ( .OUT(na2990_2), .IN1(na88_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y77     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2991_5 ( .OUT(na2991_2), .IN1(1'b0), .IN2(na99_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2992_5 ( .OUT(na2992_2), .IN1(1'b0), .IN2(na104_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2993_5 ( .OUT(na2993_2), .IN1(1'b0), .IN2(na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2994_5 ( .OUT(na2994_2), .IN1(1'b0), .IN2(na104_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2995_5 ( .OUT(na2995_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na107_2) );
// C_////Bridge      x90y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2996_5 ( .OUT(na2996_2), .IN1(na112_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2997_5 ( .OUT(na2997_2), .IN1(na121_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y64     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2998_5 ( .OUT(na2998_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na128_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2999_5 ( .OUT(na2999_2), .IN1(1'b0), .IN2(1'b0), .IN3(na129_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y108     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3000_5 ( .OUT(na3000_2), .IN1(na140_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y78     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3001_5 ( .OUT(na3001_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na152_1) );
// C_////Bridge      x80y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3002_5 ( .OUT(na3002_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na152_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3003_5 ( .OUT(na3003_2), .IN1(na176_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y83     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3004_5 ( .OUT(na3004_2), .IN1(na176_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y88     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3005_5 ( .OUT(na3005_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na176_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y66     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3006_5 ( .OUT(na3006_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na202_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y65     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3007_5 ( .OUT(na3007_2), .IN1(1'b0), .IN2(na208_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3008_5 ( .OUT(na3008_2), .IN1(1'b0), .IN2(1'b0), .IN3(na214_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3009_5 ( .OUT(na3009_2), .IN1(1'b0), .IN2(1'b0), .IN3(na214_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y99     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3010_5 ( .OUT(na3010_2), .IN1(1'b0), .IN2(1'b0), .IN3(na428_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3011_5 ( .OUT(na3011_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na429_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y82     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3012_5 ( .OUT(na3012_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na429_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3013_5 ( .OUT(na3013_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na429_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3014_5 ( .OUT(na3014_2), .IN1(1'b0), .IN2(na431_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y74     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3015_5 ( .OUT(na3015_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na433_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3016_5 ( .OUT(na3016_2), .IN1(1'b0), .IN2(na434_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y95     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3017_5 ( .OUT(na3017_2), .IN1(1'b0), .IN2(1'b0), .IN3(na438_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y78     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3018_5 ( .OUT(na3018_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na441_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3019_5 ( .OUT(na3019_2), .IN1(1'b0), .IN2(na443_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y85     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3020_5 ( .OUT(na3020_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na445_1) );
// C_////Bridge      x112y93     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3021_5 ( .OUT(na3021_2), .IN1(na448_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3022_5 ( .OUT(na3022_2), .IN1(1'b0), .IN2(1'b0), .IN3(na450_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y87     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3023_5 ( .OUT(na3023_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na450_2), .IN8(1'b0) );
// C_////Bridge      x119y97     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3024_5 ( .OUT(na3024_2), .IN1(1'b0), .IN2(1'b0), .IN3(na452_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y103     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3025_5 ( .OUT(na3025_2), .IN1(1'b0), .IN2(1'b0), .IN3(na455_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3026_5 ( .OUT(na3026_2), .IN1(1'b0), .IN2(1'b0), .IN3(na455_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3027_5 ( .OUT(na3027_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na458_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y82     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3028_5 ( .OUT(na3028_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na459_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y95     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3029_5 ( .OUT(na3029_2), .IN1(na460_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y94     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3030_5 ( .OUT(na3030_2), .IN1(1'b0), .IN2(na464_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3031_5 ( .OUT(na3031_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na472_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3032_5 ( .OUT(na3032_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na474_2) );
// C_////Bridge      x99y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3033_5 ( .OUT(na3033_2), .IN1(na475_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3034_5 ( .OUT(na3034_2), .IN1(1'b0), .IN2(na476_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3035_5 ( .OUT(na3035_2), .IN1(1'b0), .IN2(na477_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y96     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3036_5 ( .OUT(na3036_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na478_1) );
// C_////Bridge      x113y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3037_5 ( .OUT(na3037_2), .IN1(1'b0), .IN2(1'b0), .IN3(na479_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3038_5 ( .OUT(na3038_2), .IN1(1'b0), .IN2(1'b0), .IN3(na479_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3039_5 ( .OUT(na3039_2), .IN1(1'b0), .IN2(na480_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y96     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3040_5 ( .OUT(na3040_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na485_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3041_5 ( .OUT(na3041_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na489_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3042_5 ( .OUT(na3042_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na489_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3043_5 ( .OUT(na3043_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na524_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3044_5 ( .OUT(na3044_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na524_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y94     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3045_5 ( .OUT(na3045_2), .IN1(1'b0), .IN2(na527_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y81     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3046_5 ( .OUT(na3046_2), .IN1(na541_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3047_5 ( .OUT(na3047_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na544_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y85     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3048_5 ( .OUT(na3048_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na546_1) );
// C_////Bridge      x94y99     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3049_5 ( .OUT(na3049_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na557_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y105     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3050_5 ( .OUT(na3050_2), .IN1(1'b0), .IN2(na577_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3051_5 ( .OUT(na3051_2), .IN1(1'b0), .IN2(na579_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3052_5 ( .OUT(na3052_2), .IN1(1'b0), .IN2(na609_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y100     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3053_5 ( .OUT(na3053_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na621_1), .IN8(1'b0) );
// C_////Bridge      x88y104     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3054_5 ( .OUT(na3054_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na622_2), .IN8(1'b0) );
// C_////Bridge      x95y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3055_5 ( .OUT(na3055_2), .IN1(na624_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3056_5 ( .OUT(na3056_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na625_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y68     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3057_5 ( .OUT(na3057_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na626_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3058_5 ( .OUT(na3058_2), .IN1(na631_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3059_5 ( .OUT(na3059_2), .IN1(1'b0), .IN2(1'b0), .IN3(na644_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y79     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3060_5 ( .OUT(na3060_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na670_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3061_5 ( .OUT(na3061_2), .IN1(1'b0), .IN2(na686_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3062_5 ( .OUT(na3062_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na697_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3063_5 ( .OUT(na3063_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na697_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3064_5 ( .OUT(na3064_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na700_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y74     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3065_5 ( .OUT(na3065_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na700_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3066_5 ( .OUT(na3066_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na702_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3067_5 ( .OUT(na3067_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na702_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y72     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3068_5 ( .OUT(na3068_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na702_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y79     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3069_5 ( .OUT(na3069_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na702_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3070_5 ( .OUT(na3070_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na702_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3071_5 ( .OUT(na3071_2), .IN1(na703_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y69     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3072_5 ( .OUT(na3072_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na703_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y77     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3073_5 ( .OUT(na3073_2), .IN1(1'b0), .IN2(na704_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3074_5 ( .OUT(na3074_2), .IN1(1'b0), .IN2(1'b0), .IN3(na706_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3075_5 ( .OUT(na3075_2), .IN1(1'b0), .IN2(1'b0), .IN3(na709_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3076_5 ( .OUT(na3076_2), .IN1(1'b0), .IN2(na713_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3077_5 ( .OUT(na3077_2), .IN1(1'b0), .IN2(1'b0), .IN3(na719_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y68     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3078_5 ( .OUT(na3078_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na720_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3079_5 ( .OUT(na3079_2), .IN1(1'b0), .IN2(1'b0), .IN3(na724_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3080_5 ( .OUT(na3080_2), .IN1(na725_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3081_5 ( .OUT(na3081_2), .IN1(na726_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3082_5 ( .OUT(na3082_2), .IN1(na726_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3083_5 ( .OUT(na3083_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na729_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y64     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3084_5 ( .OUT(na3084_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na729_2) );
// C_////Bridge      x120y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3085_5 ( .OUT(na3085_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na735_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3086_5 ( .OUT(na3086_2), .IN1(na737_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3087_5 ( .OUT(na3087_2), .IN1(na739_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3088_5 ( .OUT(na3088_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na741_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y63     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3089_5 ( .OUT(na3089_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na743_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3090_5 ( .OUT(na3090_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na764_2), .IN8(1'b0) );
// C_////Bridge      x113y109     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3091_5 ( .OUT(na3091_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na776_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y95     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3092_5 ( .OUT(na3092_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na776_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3093_5 ( .OUT(na3093_2), .IN1(1'b0), .IN2(na779_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y98     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3094_5 ( .OUT(na3094_2), .IN1(1'b0), .IN2(na779_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y95     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3095_5 ( .OUT(na3095_2), .IN1(1'b0), .IN2(1'b0), .IN3(na780_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3096_5 ( .OUT(na3096_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na781_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y92     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3097_5 ( .OUT(na3097_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na781_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y97     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3098_5 ( .OUT(na3098_2), .IN1(1'b0), .IN2(1'b0), .IN3(na783_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y103     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3099_5 ( .OUT(na3099_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na786_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3100_5 ( .OUT(na3100_2), .IN1(1'b0), .IN2(1'b0), .IN3(na791_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y92     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3101_5 ( .OUT(na3101_2), .IN1(na800_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3102_5 ( .OUT(na3102_2), .IN1(1'b0), .IN2(na802_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y100     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3103_5 ( .OUT(na3103_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na803_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3104_5 ( .OUT(na3104_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na806_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3105_5 ( .OUT(na3105_2), .IN1(na811_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y89     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3106_5 ( .OUT(na3106_2), .IN1(1'b0), .IN2(1'b0), .IN3(na812_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3107_5 ( .OUT(na3107_2), .IN1(1'b0), .IN2(na823_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y108     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3108_5 ( .OUT(na3108_2), .IN1(na836_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y81     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3109_5 ( .OUT(na3109_2), .IN1(1'b0), .IN2(1'b0), .IN3(na850_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y101     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3110_5 ( .OUT(na3110_2), .IN1(1'b0), .IN2(1'b0), .IN3(na851_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y106     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3111_5 ( .OUT(na3111_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na853_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y107     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3112_5 ( .OUT(na3112_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na858_1) );
// C_////Bridge      x121y104     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3113_5 ( .OUT(na3113_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na858_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3114_5 ( .OUT(na3114_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na858_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y108     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3115_5 ( .OUT(na3115_2), .IN1(1'b0), .IN2(na860_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y106     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3116_5 ( .OUT(na3116_2), .IN1(1'b0), .IN2(na860_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y105     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3117_5 ( .OUT(na3117_2), .IN1(1'b0), .IN2(na863_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y110     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3118_5 ( .OUT(na3118_2), .IN1(1'b0), .IN2(na863_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y103     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3119_5 ( .OUT(na3119_2), .IN1(1'b0), .IN2(1'b0), .IN3(na877_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y106     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3120_5 ( .OUT(na3120_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na878_1), .IN8(1'b0) );
// C_////Bridge      x121y101     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3121_5 ( .OUT(na3121_2), .IN1(1'b0), .IN2(1'b0), .IN3(na878_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3122_5 ( .OUT(na3122_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na880_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y110     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3123_5 ( .OUT(na3123_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na882_1) );
// C_////Bridge      x126y110     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3124_5 ( .OUT(na3124_2), .IN1(1'b0), .IN2(na883_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y108     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3125_5 ( .OUT(na3125_2), .IN1(1'b0), .IN2(1'b0), .IN3(na884_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y103     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3126_5 ( .OUT(na3126_2), .IN1(na892_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3127_5 ( .OUT(na3127_2), .IN1(1'b0), .IN2(1'b0), .IN3(na905_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3128_5 ( .OUT(na3128_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na925_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3129_5 ( .OUT(na3129_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1010_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y94     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3130_5 ( .OUT(na3130_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1010_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y103     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3131_5 ( .OUT(na3131_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1018_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y95     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3132_5 ( .OUT(na3132_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1027_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y104     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3133_5 ( .OUT(na3133_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1031_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y83     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3134_5 ( .OUT(na3134_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1035_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3135_5 ( .OUT(na3135_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1035_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3136_5 ( .OUT(na3136_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1037_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y87     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3137_5 ( .OUT(na3137_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1039_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y81     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3138_5 ( .OUT(na3138_2), .IN1(na1045_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3139_5 ( .OUT(na3139_2), .IN1(na1045_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y87     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3140_5 ( .OUT(na3140_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1049_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3141_5 ( .OUT(na3141_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1051_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3142_5 ( .OUT(na3142_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1051_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3143_5 ( .OUT(na3143_2), .IN1(na1055_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3144_5 ( .OUT(na3144_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1065_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y107     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3145_5 ( .OUT(na3145_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1067_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y105     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3146_5 ( .OUT(na3146_2), .IN1(1'b0), .IN2(na1077_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y102     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3147_5 ( .OUT(na3147_2), .IN1(1'b0), .IN2(na1077_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y107     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3148_5 ( .OUT(na3148_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1081_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y102     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3149_5 ( .OUT(na3149_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1081_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y110     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3150_5 ( .OUT(na3150_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1083_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y95     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3151_5 ( .OUT(na3151_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1083_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y105     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3152_5 ( .OUT(na3152_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1084_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y106     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3153_5 ( .OUT(na3153_2), .IN1(na1085_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3154_5 ( .OUT(na3154_2), .IN1(na1087_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y79     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3155_5 ( .OUT(na3155_2), .IN1(na1087_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3156_5 ( .OUT(na3156_2), .IN1(na1087_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3157_5 ( .OUT(na3157_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1089_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3158_5 ( .OUT(na3158_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1089_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3159_5 ( .OUT(na3159_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1099_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3160_5 ( .OUT(na3160_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1103_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y106     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3161_5 ( .OUT(na3161_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1270_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y70     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3162_5 ( .OUT(na3162_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1273_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y70     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3163_5 ( .OUT(na3163_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1458_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y100     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3164_5 ( .OUT(na3164_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1461_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y108     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3165_5 ( .OUT(na3165_2), .IN1(na1465_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y109     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3166_5 ( .OUT(na3166_2), .IN1(na1465_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3167_5 ( .OUT(na3167_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2407_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y93     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3168_5 ( .OUT(na3168_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2409_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y107     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3169_5 ( .OUT(na3169_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2410_1) );
// C_////Bridge      x81y95     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3170_5 ( .OUT(na3170_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2410_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y88     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3171_5 ( .OUT(na3171_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2410_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y102     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3172_5 ( .OUT(na3172_2), .IN1(1'b0), .IN2(na2413_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y77     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3173_5 ( .OUT(na3173_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2414_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3174_5 ( .OUT(na3174_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2416_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3175_5 ( .OUT(na3175_2), .IN1(na2423_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y75     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3176_5 ( .OUT(na3176_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2426_1) );
// C_////Bridge      x80y85     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3177_5 ( .OUT(na3177_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2446_1) );
// C_////Bridge      x87y78     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3178_5 ( .OUT(na3178_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2474_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y97     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3179_5 ( .OUT(na3179_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2518_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y85     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3180_5 ( .OUT(na3180_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2529_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y89     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3181_5 ( .OUT(na3181_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2549_1) );
// C_////Bridge      x93y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3182_5 ( .OUT(na3182_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2565_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y109     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3183_5 ( .OUT(na3183_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2629_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y67     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3184_5 ( .OUT(na3184_2), .IN1(na2680_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y82     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3185_5 ( .OUT(na3185_2), .IN1(na2691_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y68     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3186_5 ( .OUT(na3186_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2693_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y63     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3187_5 ( .OUT(na3187_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2694_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y64     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3188_5 ( .OUT(na3188_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2694_2), .IN8(1'b0) );
// C_////Bridge      x107y92     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3189_5 ( .OUT(na3189_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2697_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y80     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3190_5 ( .OUT(na3190_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2698_2), .IN8(1'b0) );
// C_////Bridge      x103y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3191_5 ( .OUT(na3191_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2701_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3192_5 ( .OUT(na3192_2), .IN1(na2702_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3193_5 ( .OUT(na3193_2), .IN1(na2703_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3194_5 ( .OUT(na3194_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2704_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3195_5 ( .OUT(na3195_2), .IN1(na2705_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y101     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3196_5 ( .OUT(na3196_2), .IN1(na2707_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3197_5 ( .OUT(na3197_2), .IN1(na2718_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y95     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3198_5 ( .OUT(na3198_2), .IN1(na2718_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3199_5 ( .OUT(na3199_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2729_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y108     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3200_5 ( .OUT(na3200_2), .IN1(na2746_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y105     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3201_5 ( .OUT(na3201_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2751_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y108     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3202_5 ( .OUT(na3202_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2757_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y108     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3203_5 ( .OUT(na3203_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2757_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y106     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3204_5 ( .OUT(na3204_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2758_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3205_5 ( .OUT(na3205_2), .IN1(na2763_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y98     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3206_5 ( .OUT(na3206_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2771_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y105     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3207_5 ( .OUT(na3207_2), .IN1(1'b0), .IN2(na2774_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y104     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3208_5 ( .OUT(na3208_2), .IN1(na2775_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y92     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3209_5 ( .OUT(na3209_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2778_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3210_5 ( .OUT(na3210_2), .IN1(na2779_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3211_5 ( .OUT(na3211_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2780_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3212_5 ( .OUT(na3212_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2781_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3213_5 ( .OUT(na3213_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2782_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3214_5 ( .OUT(na3214_2), .IN1(1'b0), .IN2(na2855_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y107     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3215_5 ( .OUT(na3215_2), .IN1(1'b0), .IN2(na2908_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3216_5 ( .OUT(na3216_2), .IN1(1'b0), .IN2(na2923_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y80     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3217_5 ( .OUT(na3217_2), .IN1(1'b0), .IN2(na2923_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y100     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a3218_5 ( .OUT(na3218_2), .IN1(na2930_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_CP_route////      x80y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3219_1 ( .OUT(na3219_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x81y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3220_1 ( .OUT(na3220_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x82y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3221_1 ( .OUT(na3221_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x83y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3222_1 ( .OUT(na3222_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x84y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3223_1 ( .OUT(na3223_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x85y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3224_1 ( .OUT(na3224_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x86y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3225_1 ( .OUT(na3225_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x87y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3226_1 ( .OUT(na3226_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x88y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3227_1 ( .OUT(na3227_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x89y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3228_1 ( .OUT(na3228_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x90y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3229_1 ( .OUT(na3229_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x91y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3230_1 ( .OUT(na3230_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x92y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3231_1 ( .OUT(na3231_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x93y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3232_1 ( .OUT(na3232_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x94y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3233_1 ( .OUT(na3233_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x95y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3234_1 ( .OUT(na3234_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x96y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3235_1 ( .OUT(na3235_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x97y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3236_1 ( .OUT(na3236_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x98y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3237_1 ( .OUT(na3237_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x99y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3238_1 ( .OUT(na3238_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x100y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3239_1 ( .OUT(na3239_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x101y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3240_1 ( .OUT(na3240_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x102y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3241_1 ( .OUT(na3241_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x103y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3242_1 ( .OUT(na3242_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x104y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3243_1 ( .OUT(na3243_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x105y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3244_1 ( .OUT(na3244_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x106y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3245_1 ( .OUT(na3245_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x107y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3246_1 ( .OUT(na3246_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x108y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3247_1 ( .OUT(na3247_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x109y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3248_1 ( .OUT(na3248_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x110y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3249_1 ( .OUT(na3249_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x111y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3250_1 ( .OUT(na3250_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x112y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3251_1 ( .OUT(na3251_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x113y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3252_1 ( .OUT(na3252_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x114y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3253_1 ( .OUT(na3253_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x115y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3254_1 ( .OUT(na3254_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x116y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3255_1 ( .OUT(na3255_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x117y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3256_1 ( .OUT(na3256_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x118y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3257_1 ( .OUT(na3257_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x119y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3258_1 ( .OUT(na3258_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x120y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3259_1 ( .OUT(na3259_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x121y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3260_1 ( .OUT(na3260_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x122y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3261_1 ( .OUT(na3261_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_CP_route////      x123y60     80'h00_0018_24_7000_0C00_0000
C_CP_route #(.CPE_CFG (9'b0_0000_0000)) 
           _a3262_1 ( .OUT(na3262_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x79y60     80'h00_0078_09_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3263_1 ( .OUT(na3263_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1487_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3263_4 ( .OUT(na3263_2), .IN1(1'b1), .IN2(na62_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9000)) 
           _a3263_6 ( .COUTX(na3263_3), .POUTX(na3263_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na3263_1), .OUT2(na3263_2), .COMP_OUT(1'b0) );
endmodule
